`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: TEC
// Engineer: Steven Astorga - Steven Avila - Luis Saborio
// Module Name: Memoria simulada para pruebas varias
//////////////////////////////////////////////////////////////////////////////////
module memoria(
			input clk,
			input wire [10:0] dir,
			output reg [31:0] dato
);
reg [10:0] addr_reg; 
   // body
   always @(posedge clk) 
      addr_reg <= dir;

	always @*
      case (addr_reg)
			11'h0 : dato = 32'b11111111111111111111111111111111;
			11'h1 : dato = 32'b11111111111111111111111111111111;
			11'h2 : dato = 32'b11111111111111111111111111111111;
			11'h3 : dato = 32'b11111111111111111111111111111111;
			11'h4 : dato = 32'b11111111111111111111111111111111;
			11'h5 : dato = 32'b11111111111111111111111111111111;
			11'h6 : dato = 32'b11111111111111111111111111111111;
			11'h7 : dato = 32'b11111111111111111111111111111111;
			11'h8 : dato = 32'b11111111111111111111111111111111;
			11'h9 : dato = 32'b11111111111111111111111111111111;
			11'ha : dato = 32'b11111111111111111111111111111111;
			11'hb : dato = 32'b11111111111111111111111111111111;
			11'hc : dato = 32'b11111111111111111111111111111111;
			11'hd : dato = 32'b11111111111111111111111111111111;
			11'he : dato = 32'b11111111111111111111111111111111;
			11'hf : dato = 32'b11111111111111111111111111111111;
			11'h10 : dato = 32'b11111111111111111111111111111111;
			11'h11 : dato = 32'b11111111111111111111111111111111;
			11'h12 : dato = 32'b11111111111111111111111111111111;
			11'h13 : dato = 32'b11111111111111111111111111111111;
			11'h14 : dato = 32'b11111111111111111111111111111111;
			11'h15 : dato = 32'b11111111111111111111111111111111;
			11'h16 : dato = 32'b11111111111111111111111111111111;
			11'h17 : dato = 32'b11111111111111111111111111111111;
			11'h18 : dato = 32'b11111111111111111111111111111111;
			11'h19 : dato = 32'b11111111111111111111111111111111;
			11'h1a : dato = 32'b11111111111111111111111111111111;
			11'h1b : dato = 32'b11111111111111111111111111111111;
			11'h1c : dato = 32'b11111111111111111111111111111111;
			11'h1d : dato = 32'b11111111111111111111111111111111;
			11'h1e : dato = 32'b11111111111111111111111111111111;
			11'h1f : dato = 32'b11111111111111111111111111111111;
			11'h20 : dato = 32'b11111111111111111111111111111111;
			11'h21 : dato = 32'b11111111111111111111111111111111;
			11'h22 : dato = 32'b11111111111111111111111111111111;
			11'h23 : dato = 32'b11111111111111111111111111111111;
			11'h24 : dato = 32'b11111111111111111111111111111111;
			11'h25 : dato = 32'b11111111111111111111111111111111;
			11'h26 : dato = 32'b11111111111111111111111111111111;
			11'h27 : dato = 32'b11111111111111111111111111111111;
			11'h28 : dato = 32'b11111111111111111111111111111111;
			11'h29 : dato = 32'b11111111111111111111111111111111;
			11'h2a : dato = 32'b11111111111111111111111111111111;
			11'h2b : dato = 32'b11111111111111111111111111111111;
			11'h2c : dato = 32'b11111111111111111111111111111111;
			11'h2d : dato = 32'b11111111111111111111111111111111;
			11'h2e : dato = 32'b11111111111111111111111111111111;
			11'h2f : dato = 32'b11111111111111111111111111111111;
			11'h30 : dato = 32'b11111111111111111111111111111111;
			11'h31 : dato = 32'b11111111111111111111111111111111;
			11'h32 : dato = 32'b11111111111111111111111111111111;
			11'h33 : dato = 32'b11111111111111111111111111111111;
			11'h34 : dato = 32'b11111111111111111110111110111110;
			11'h35 : dato = 32'b10011000011111001100110111111111;
			11'h36 : dato = 32'b11111111111111111111111111111111;
			11'h37 : dato = 32'b11111111111111111111111111111111;
			11'h38 : dato = 32'b11111111111111111111111111111111;
			11'h39 : dato = 32'b11111111111111111111111111111111;
			11'h3a : dato = 32'b11111111111111111111111111111111;
			11'h3b : dato = 32'b11111111111111111111111111111111;
			11'h3c : dato = 32'b11111111111111111111111111111111;
			11'h3d : dato = 32'b11111111111111111111111111111111;
			11'h3e : dato = 32'b11111111111111111111111111111111;
			11'h3f : dato = 32'b11111111111111111111111111111111;
			11'h40 : dato = 32'b11111111111111111111111111111111;
			11'h41 : dato = 32'b11111111111111111111111111111111;
			11'h42 : dato = 32'b11111111111111111111111111111111;
			11'h43 : dato = 32'b11111111111111111111111111111111;
			11'h44 : dato = 32'b11111111111111111111111111111111;
			11'h45 : dato = 32'b11111111111111111111111111111111;
			11'h46 : dato = 32'b11111111111111111111111111111111;
			11'h47 : dato = 32'b11111111111111111111111111111111;
			11'h48 : dato = 32'b11011111100101100110100001100110;
			11'h49 : dato = 32'b01100110011001101100100011111111;
			11'h4a : dato = 32'b11111111111111111111111111111111;
			11'h4b : dato = 32'b11111111111111111111111111111111;
			11'h4c : dato = 32'b11111111111111111111111111111111;
			11'h4d : dato = 32'b11111111111111111111111111111111;
			11'h4e : dato = 32'b11111111111111111111111111111111;
			11'h4f : dato = 32'b11111111111111111111111111111111;
			11'h50 : dato = 32'b11111111111111111111111111111111;
			11'h51 : dato = 32'b11111111111111111111111111111111;
			11'h52 : dato = 32'b11111111111111111111111111111111;
			11'h53 : dato = 32'b11111111111111111111111111111111;
			11'h54 : dato = 32'b11111111111111111111111111111111;
			11'h55 : dato = 32'b11111111111111111111111111111111;
			11'h56 : dato = 32'b11111111111111111111111111111111;
			11'h57 : dato = 32'b11111111111111111111111111111111;
			11'h58 : dato = 32'b11111111111111111111111111111111;
			11'h59 : dato = 32'b11111111111111111111111111111111;
			11'h5a : dato = 32'b11111111111111111111111111111111;
			11'h5b : dato = 32'b11111111111111111111001010011111;
			11'h5c : dato = 32'b01100110011001100110011001100110;
			11'h5d : dato = 32'b01100110011001101100111011111111;
			11'h5e : dato = 32'b11111111111111111111111111111111;
			11'h5f : dato = 32'b11111111111111111111111111111111;
			11'h60 : dato = 32'b11111111111111111111111111111111;
			11'h61 : dato = 32'b11111111111111111111111111111111;
			11'h62 : dato = 32'b11111111111111111111111111111111;
			11'h63 : dato = 32'b11111111111111111111111111111111;
			11'h64 : dato = 32'b11111111111111111111111111111111;
			11'h65 : dato = 32'b11111111111111111111111111111111;
			11'h66 : dato = 32'b11111111111111111111111111111111;
			11'h67 : dato = 32'b11111111111111111111111111111111;
			11'h68 : dato = 32'b11111111111111111111111111111111;
			11'h69 : dato = 32'b11111111111111111111111111111111;
			11'h6a : dato = 32'b11111111111111111111111111111111;
			11'h6b : dato = 32'b11111111111111111111111111111111;
			11'h6c : dato = 32'b11111111111111111111111111111111;
			11'h6d : dato = 32'b11111111111111111111111111111111;
			11'h6e : dato = 32'b11111111111111111111111111111111;
			11'h6f : dato = 32'b11111111110011010110111001100110;
			11'h70 : dato = 32'b01100110011001100110011001100110;
			11'h71 : dato = 32'b01100110011001101101101011111111;
			11'h72 : dato = 32'b11111111111111111111111111111111;
			11'h73 : dato = 32'b11111111111111111111111111111111;
			11'h74 : dato = 32'b11111111111111111111111111111111;
			11'h75 : dato = 32'b11111111111111111111111111111111;
			11'h76 : dato = 32'b11111111111111111111111111111111;
			11'h77 : dato = 32'b11111111111111111111111111111111;
			11'h78 : dato = 32'b11111111111111111111111111111111;
			11'h79 : dato = 32'b11111111111111111111111111111111;
			11'h7a : dato = 32'b11111111111111111111111111111111;
			11'h7b : dato = 32'b11111111111111111111111111111111;
			11'h7c : dato = 32'b11111111111111111111111111111111;
			11'h7d : dato = 32'b11111111111111111111111111111111;
			11'h7e : dato = 32'b11111111111111111111111111111111;
			11'h7f : dato = 32'b11111111111111111111111111111111;
			11'h80 : dato = 32'b11111111111111111111111111111111;
			11'h81 : dato = 32'b11111111111111111111111111111111;
			11'h82 : dato = 32'b11111111111111111111111111111111;
			11'h83 : dato = 32'b11010101011001110110011001100110;
			11'h84 : dato = 32'b01100110011001100110011001100110;
			11'h85 : dato = 32'b01100110011001101110111111111111;
			11'h86 : dato = 32'b11111111111111111111111111111111;
			11'h87 : dato = 32'b11111111111111111111111111111111;
			11'h88 : dato = 32'b11111111111111111111111111111111;
			11'h89 : dato = 32'b11111111111111111111111111111111;
			11'h8a : dato = 32'b11111111111111111111111111111111;
			11'h8b : dato = 32'b11111111111111111111111111111111;
			11'h8c : dato = 32'b11111111111111111111111111111111;
			11'h8d : dato = 32'b11111111111111111111111111111111;
			11'h8e : dato = 32'b11111111111111111111111111111111;
			11'h8f : dato = 32'b11111111111111111111111111111111;
			11'h90 : dato = 32'b11111111111111111111111111111111;
			11'h91 : dato = 32'b11111111111111111111111111111111;
			11'h92 : dato = 32'b11111111111111111111111111111111;
			11'h93 : dato = 32'b11111111111111111111111111111111;
			11'h94 : dato = 32'b11111111111111111111111111111111;
			11'h95 : dato = 32'b11111111111111111111111111111111;
			11'h96 : dato = 32'b11111111111111111111111111100110;
			11'h97 : dato = 32'b01110000011001100110011001100110;
			11'h98 : dato = 32'b01100110011001100110011001100110;
			11'h99 : dato = 32'b01100110011100101111111111111111;
			11'h9a : dato = 32'b11111111111111111111111111111111;
			11'h9b : dato = 32'b11111111111111111111111111111111;
			11'h9c : dato = 32'b11111111111111111111111111111111;
			11'h9d : dato = 32'b11111111111111111111111111111111;
			11'h9e : dato = 32'b11111111111111111111111111111111;
			11'h9f : dato = 32'b11111111111111111111111111111111;
			11'ha0 : dato = 32'b11111111111111111111111111111111;
			11'ha1 : dato = 32'b11111111111111111111111111111111;
			11'ha2 : dato = 32'b11111111111111111111111111111111;
			11'ha3 : dato = 32'b11111111111111111111111111111111;
			11'ha4 : dato = 32'b11111111111111111111111111111111;
			11'ha5 : dato = 32'b11111111111111111111111111111111;
			11'ha6 : dato = 32'b11111111111111111111111111111111;
			11'ha7 : dato = 32'b11111111111111111111111111111111;
			11'ha8 : dato = 32'b11111111111111111111111111111111;
			11'ha9 : dato = 32'b11111111111111111111111111111111;
			11'haa : dato = 32'b11111111111111111110110101111001;
			11'hab : dato = 32'b01100110011001100110011001100110;
			11'hac : dato = 32'b01100110011001100110011001100110;
			11'had : dato = 32'b01100110100111101111111111111111;
			11'hae : dato = 32'b11111111111111111111111111111111;
			11'haf : dato = 32'b11111111111111111111111111111111;
			11'hb0 : dato = 32'b11111111111111111111111111111111;
			11'hb1 : dato = 32'b11111111111111111111111111111111;
			11'hb2 : dato = 32'b11111111111111111111111111111111;
			11'hb3 : dato = 32'b11111111111111111111111111111111;
			11'hb4 : dato = 32'b11111111111111111111111111111111;
			11'hb5 : dato = 32'b11111111111111111111111111111111;
			11'hb6 : dato = 32'b11111111111111111111111111111111;
			11'hb7 : dato = 32'b11111111111111111111111111111111;
			11'hb8 : dato = 32'b11111111111111111111111111111111;
			11'hb9 : dato = 32'b11111111111111111111111111111111;
			11'hba : dato = 32'b11111111111111111111111111111111;
			11'hbb : dato = 32'b11111111111111111111111111111111;
			11'hbc : dato = 32'b11111111111111111111111111111111;
			11'hbd : dato = 32'b11111111111111111111111111111111;
			11'hbe : dato = 32'b11111111111100110111101101100110;
			11'hbf : dato = 32'b01100110011001100110011001100110;
			11'hc0 : dato = 32'b01100110011001100110011001100110;
			11'hc1 : dato = 32'b01100110110101111111111111111111;
			11'hc2 : dato = 32'b11111111111111111111111111111111;
			11'hc3 : dato = 32'b11111111111111111111111111111111;
			11'hc4 : dato = 32'b11111111111111111111111111111111;
			11'hc5 : dato = 32'b11111111111111111111111111111111;
			11'hc6 : dato = 32'b11111111111111111111111111111111;
			11'hc7 : dato = 32'b11111111111111111111111111111111;
			11'hc8 : dato = 32'b11111111111111111111111111111111;
			11'hc9 : dato = 32'b11111111111111111111111111111111;
			11'hca : dato = 32'b11111111111111111111111111111111;
			11'hcb : dato = 32'b11111111111111111111111111111111;
			11'hcc : dato = 32'b11111111111111111111111111111111;
			11'hcd : dato = 32'b11111111111111111111111111111111;
			11'hce : dato = 32'b11111111111111111111111111111111;
			11'hcf : dato = 32'b11111111111111111111111111111111;
			11'hd0 : dato = 32'b11111111111111111111111111111111;
			11'hd1 : dato = 32'b11111111111111111111111111111111;
			11'hd2 : dato = 32'b11111111100111100110011001100110;
			11'hd3 : dato = 32'b01100110011001100110011001100110;
			11'hd4 : dato = 32'b01100110011001100110011001100110;
			11'hd5 : dato = 32'b10000011111111111111111111111111;
			11'hd6 : dato = 32'b11111111111111111111111111111111;
			11'hd7 : dato = 32'b11111111111111111111111111111111;
			11'hd8 : dato = 32'b11111111111111111111111111111111;
			11'hd9 : dato = 32'b11111111111111111111111111111111;
			11'hda : dato = 32'b11111111111111111111111111111111;
			11'hdb : dato = 32'b11111111111111111111111111111111;
			11'hdc : dato = 32'b11111111111111111111111111111111;
			11'hdd : dato = 32'b11111111111111111111111111111111;
			11'hde : dato = 32'b11111111111111111111111111111111;
			11'hdf : dato = 32'b11111111111111111111111111111111;
			11'he0 : dato = 32'b11111111111111111111111111111111;
			11'he1 : dato = 32'b11111111111111111111111111111111;
			11'he2 : dato = 32'b11111111111111111111111111111111;
			11'he3 : dato = 32'b11111111111111111111111111111111;
			11'he4 : dato = 32'b11111111111111111111111111111111;
			11'he5 : dato = 32'b11111111111111111111111111111111;
			11'he6 : dato = 32'b11101001011001110110011001100110;
			11'he7 : dato = 32'b01100110011001100110011001100110;
			11'he8 : dato = 32'b01100110011001100110011001100110;
			11'he9 : dato = 32'b11001001111111111111111111111111;
			11'hea : dato = 32'b11111111111111111111111111111111;
			11'heb : dato = 32'b11111111111111111111111111111111;
			11'hec : dato = 32'b11111111111111111111111111111111;
			11'hed : dato = 32'b11111111111111111111111111111111;
			11'hee : dato = 32'b11111111111111111111111111111111;
			11'hef : dato = 32'b11111111111111111111111111111111;
			11'hf0 : dato = 32'b11111111111111111111111111111111;
			11'hf1 : dato = 32'b11111111111111111111111111111111;
			11'hf2 : dato = 32'b11111111111111111111111111111111;
			11'hf3 : dato = 32'b11111111111111111111111111111111;
			11'hf4 : dato = 32'b11111111111111111111111111111111;
			11'hf5 : dato = 32'b11111111111111111111111111111111;
			11'hf6 : dato = 32'b11111111111111111111111111111111;
			11'hf7 : dato = 32'b11111111111111111111111111111111;
			11'hf8 : dato = 32'b11111111111111111111111111111111;
			11'hf9 : dato = 32'b11111111111111111111111111111111;
			11'hfa : dato = 32'b10101010011001100110011001100110;
			11'hfb : dato = 32'b01100110011001100110011001100110;
			11'hfc : dato = 32'b01100110011001100110011010001111;
			11'hfd : dato = 32'b11111101111111111111111111111111;
			11'hfe : dato = 32'b11111111111111111111111111111111;
			11'hff : dato = 32'b11111111111111111111111111111111;
			11'h100 : dato = 32'b11111111111111111111111111111111;
			11'h101 : dato = 32'b11111111111111111111111111111111;
			11'h102 : dato = 32'b11111111111111111111111111111111;
			11'h103 : dato = 32'b11111111111111111111111111111111;
			11'h104 : dato = 32'b11111111111111111111111111111111;
			11'h105 : dato = 32'b11111111111111111111111111111111;
			11'h106 : dato = 32'b11111111111111111111111111111111;
			11'h107 : dato = 32'b11111111111111111111111111111111;
			11'h108 : dato = 32'b11111111111111111111111111111111;
			11'h109 : dato = 32'b11111111111111111111111111111111;
			11'h10a : dato = 32'b11111111111111111111111111111111;
			11'h10b : dato = 32'b11111111111111111111111111111111;
			11'h10c : dato = 32'b11111111111111111111111111111111;
			11'h10d : dato = 32'b11111111111111111111111111111100;
			11'h10e : dato = 32'b01110001011001100110011001100110;
			11'h10f : dato = 32'b01100110011001100110011001100110;
			11'h110 : dato = 32'b01100110011001101000001011111001;
			11'h111 : dato = 32'b11111111111111111111111111111111;
			11'h112 : dato = 32'b11111111111111111111111111111111;
			11'h113 : dato = 32'b11111111111111111111111111111111;
			11'h114 : dato = 32'b11111111111111111111111111111111;
			11'h115 : dato = 32'b11111111111111111111111111111111;
			11'h116 : dato = 32'b11111111111111111111111111111111;
			11'h117 : dato = 32'b11111111111111111111111111111111;
			11'h118 : dato = 32'b11111111111111111111111111111111;
			11'h119 : dato = 32'b11111111111111111111111111111111;
			11'h11a : dato = 32'b11111111111111111111111111111111;
			11'h11b : dato = 32'b11111111111111111111111111111111;
			11'h11c : dato = 32'b11111111111111111111111111111111;
			11'h11d : dato = 32'b11111111111111111111111111111111;
			11'h11e : dato = 32'b11111111111111111111111111111111;
			11'h11f : dato = 32'b11111111111111111111111111111111;
			11'h120 : dato = 32'b11111111111111111111111111111111;
			11'h121 : dato = 32'b11111111111111111111111111011010;
			11'h122 : dato = 32'b01100110011001100110011001100110;
			11'h123 : dato = 32'b01100110011001100110011001100110;
			11'h124 : dato = 32'b01100110011101001110110011111111;
			11'h125 : dato = 32'b11111111111111111111111111111111;
			11'h126 : dato = 32'b11111111111111111111111111111111;
			11'h127 : dato = 32'b11111111111111111111111111111111;
			11'h128 : dato = 32'b11111111111111111111111111111111;
			11'h129 : dato = 32'b11111111111111111111111111111111;
			11'h12a : dato = 32'b11111111111111111111111111111111;
			11'h12b : dato = 32'b11111111111111111111111111111111;
			11'h12c : dato = 32'b11111111111111111111111111111111;
			11'h12d : dato = 32'b11111111111111111111111111111111;
			11'h12e : dato = 32'b11111111111111111111111111111111;
			11'h12f : dato = 32'b11111111111111111111111111111111;
			11'h130 : dato = 32'b11111111111111111111111111111111;
			11'h131 : dato = 32'b11111111111111111111111111111111;
			11'h132 : dato = 32'b11111111111111111111111111111111;
			11'h133 : dato = 32'b11111111111111111111111111111111;
			11'h134 : dato = 32'b11111111111111111111111111111111;
			11'h135 : dato = 32'b11111111111111111111111110111100;
			11'h136 : dato = 32'b01100110011001100110011001100110;
			11'h137 : dato = 32'b01100110011001100110011001100110;
			11'h138 : dato = 32'b01100111110110001111111111111111;
			11'h139 : dato = 32'b11111111111111111111111111111111;
			11'h13a : dato = 32'b11111111111111111111111111111111;
			11'h13b : dato = 32'b11111111111111111111111111111111;
			11'h13c : dato = 32'b11111111111111111111111111111111;
			11'h13d : dato = 32'b11111111111111111111111111111111;
			11'h13e : dato = 32'b11111111111111111111111111111111;
			11'h13f : dato = 32'b11111111111111111111111111111111;
			11'h140 : dato = 32'b11111111111111111111111111111111;
			11'h141 : dato = 32'b11111111111111111111111111111111;
			11'h142 : dato = 32'b11111111111111111111111111111111;
			11'h143 : dato = 32'b11111111111111111111111111111111;
			11'h144 : dato = 32'b11111111111111111111111111111111;
			11'h145 : dato = 32'b11111111111111111111111111111111;
			11'h146 : dato = 32'b11111111111111111111111111111111;
			11'h147 : dato = 32'b11111111111111111111111111111111;
			11'h148 : dato = 32'b11111111111111111111111111111111;
			11'h149 : dato = 32'b11111111111111111111111110101001;
			11'h14a : dato = 32'b01100110011001100110011001100110;
			11'h14b : dato = 32'b01100110011001100110011001101100;
			11'h14c : dato = 32'b11001100111111111111111111111111;
			11'h14d : dato = 32'b11111111111111111111111111111111;
			11'h14e : dato = 32'b11111111111111111111111111111111;
			11'h14f : dato = 32'b11111111111111111111111111111111;
			11'h150 : dato = 32'b11111111111111111111111111111111;
			11'h151 : dato = 32'b11111111111111111111111111111111;
			11'h152 : dato = 32'b11111111111111111111111111111111;
			11'h153 : dato = 32'b11111111111111111111111111111111;
			11'h154 : dato = 32'b11111111111111111111111111111111;
			11'h155 : dato = 32'b11111111111111111111111111111111;
			11'h156 : dato = 32'b11111111111111111111111111111111;
			11'h157 : dato = 32'b11111111111111111111111111111111;
			11'h158 : dato = 32'b11111111111111111111111111111111;
			11'h159 : dato = 32'b11111111111111111111111111111111;
			11'h15a : dato = 32'b11111111111111111111111111111111;
			11'h15b : dato = 32'b11111111111111111111111111111111;
			11'h15c : dato = 32'b11111111111111111111111111111111;
			11'h15d : dato = 32'b11111111111111111111111110100001;
			11'h15e : dato = 32'b01100110011001100110011001100110;
			11'h15f : dato = 32'b01100110011001101000110011100011;
			11'h160 : dato = 32'b11111111111111111111111111111111;
			11'h161 : dato = 32'b11111111111111111111111111111111;
			11'h162 : dato = 32'b11111111111111111111111111111111;
			11'h163 : dato = 32'b11111111111111111111111111111111;
			11'h164 : dato = 32'b11111111111111111111111111111111;
			11'h165 : dato = 32'b11111111111111111111111111111111;
			11'h166 : dato = 32'b11111111111111111111111111111111;
			11'h167 : dato = 32'b11111111111111111111111111111111;
			11'h168 : dato = 32'b11111111111111111111111111111111;
			11'h169 : dato = 32'b11111111111111111111111111111111;
			11'h16a : dato = 32'b11111111111111111111111111111111;
			11'h16b : dato = 32'b11111111111111111111111111111111;
			11'h16c : dato = 32'b11111111111111111111111111111111;
			11'h16d : dato = 32'b11111111111111111111111111111111;
			11'h16e : dato = 32'b11111111111111111111111111111111;
			11'h16f : dato = 32'b11111111111111111111111111111111;
			11'h170 : dato = 32'b11111111111111111111111111111111;
			11'h171 : dato = 32'b11111111111111111111111110100010;
			11'h172 : dato = 32'b01100110011001100110011001101010;
			11'h173 : dato = 32'b10010101110110111111111111111111;
			11'h174 : dato = 32'b11111111111111111111111111111111;
			11'h175 : dato = 32'b11111111111111111111111111111111;
			11'h176 : dato = 32'b11111111111111111111111111111111;
			11'h177 : dato = 32'b11111111111111111111111111111111;
			11'h178 : dato = 32'b11111111111111111111111111111111;
			11'h179 : dato = 32'b11111111111111111111111111111111;
			11'h17a : dato = 32'b11111111111111111111111111111111;
			11'h17b : dato = 32'b11111111111111111111111111111111;
			11'h17c : dato = 32'b11111111111111111111111111111111;
			11'h17d : dato = 32'b11111111111111111111111111111111;
			11'h17e : dato = 32'b11111111111111111111111111111111;
			11'h17f : dato = 32'b11111111111111111111111111111111;
			11'h180 : dato = 32'b11111111111111111111111111111111;
			11'h181 : dato = 32'b11111111111111111111111111111111;
			11'h182 : dato = 32'b11111111111111111111111111111111;
			11'h183 : dato = 32'b11111111111111111111111111111111;
			11'h184 : dato = 32'b11111111111111111111111111111111;
			11'h185 : dato = 32'b11111111111111111111111111011100;
			11'h186 : dato = 32'b10110110101110011100111111110101;
			11'h187 : dato = 32'b11111111111111111111111111111111;
			11'h188 : dato = 32'b11111111111111111111111111111111;
			11'h189 : dato = 32'b11111111111111111111111111111111;
			11'h18a : dato = 32'b11111111111111111111111111111111;
			11'h18b : dato = 32'b11111111111111111111111111111111;
			11'h18c : dato = 32'b11111111111111111111111111111111;
			11'h18d : dato = 32'b11111111111111111111111111111111;
			11'h18e : dato = 32'b11111111111111111111111111111111;
			11'h18f : dato = 32'b11111111111111111111111111111111;
			11'h190 : dato = 32'b11111111111111111111111111111111;
			11'h191 : dato = 32'b11111111111111111111111111111111;
			11'h192 : dato = 32'b11111111111111111111111111111111;
			11'h193 : dato = 32'b11111111111111111111111111111111;
			11'h194 : dato = 32'b11111111111111111111111111111111;
			11'h195 : dato = 32'b11111111111111111111111111100011;
			11'h196 : dato = 32'b10111110101000111001000010001001;
			11'h197 : dato = 32'b10001111101001101100111111111010;
			11'h198 : dato = 32'b11111111111111111111111111111111;
			11'h199 : dato = 32'b11111111111111111111111111111111;
			11'h19a : dato = 32'b11111111111111111111111111111111;
			11'h19b : dato = 32'b11111111111111111111111111111111;
			11'h19c : dato = 32'b11100111101110011001001001111011;
			11'h19d : dato = 32'b01101000011001100110011101111000;
			11'h19e : dato = 32'b10001100101100001101111111111111;
			11'h19f : dato = 32'b11111111111111111111111111111111;
			11'h1a0 : dato = 32'b11111111111111111111111111111111;
			11'h1a1 : dato = 32'b11111111111111111111111111111111;
			11'h1a2 : dato = 32'b11111111111111111111111111111111;
			11'h1a3 : dato = 32'b11111111111111111111111111111111;
			11'h1a4 : dato = 32'b11111111111111111111111111111111;
			11'h1a5 : dato = 32'b11111111111111111111111111111111;
			11'h1a6 : dato = 32'b11111111111111111111111111111111;
			11'h1a7 : dato = 32'b11111111111111111111111111111111;
			11'h1a8 : dato = 32'b11111111111111111111111111111111;
			11'h1a9 : dato = 32'b11101001101100100111101101100110;
			11'h1aa : dato = 32'b01100110011001100110011001100110;
			11'h1ab : dato = 32'b01100110011001100110011001101100;
			11'h1ac : dato = 32'b10010100101111001110100111111111;
			11'h1ad : dato = 32'b11111111111111111111111111111111;
			11'h1ae : dato = 32'b11111111111111111111111111111111;
			11'h1af : dato = 32'b11111001110011001010001001111011;
			11'h1b0 : dato = 32'b01100110011001100110011001100110;
			11'h1b1 : dato = 32'b01100110011001100110011001100110;
			11'h1b2 : dato = 32'b01100110011001100110011001110110;
			11'h1b3 : dato = 32'b10100111111010001111111111111111;
			11'h1b4 : dato = 32'b11111111111111111111111111111111;
			11'h1b5 : dato = 32'b11111111111111111111111111111111;
			11'h1b6 : dato = 32'b11111111111111111111111111111111;
			11'h1b7 : dato = 32'b11111111111111111111111111111111;
			11'h1b8 : dato = 32'b11111111111111111111111111111111;
			11'h1b9 : dato = 32'b11111111111111111111111111111111;
			11'h1ba : dato = 32'b11111111111111111111111111111111;
			11'h1bb : dato = 32'b11111111111111111111111111111111;
			11'h1bc : dato = 32'b11111111111111111110101110011111;
			11'h1bd : dato = 32'b01100110011001100110011001100110;
			11'h1be : dato = 32'b01100110011001100110011001100110;
			11'h1bf : dato = 32'b01100110011001100110011001100110;
			11'h1c0 : dato = 32'b01100110011001100110011010000011;
			11'h1c1 : dato = 32'b10110110111000101111111011111111;
			11'h1c2 : dato = 32'b11111111111110111101000110011110;
			11'h1c3 : dato = 32'b01101101011001100110011001100110;
			11'h1c4 : dato = 32'b01100110011001100110011001100110;
			11'h1c5 : dato = 32'b01100110011001100110011001100110;
			11'h1c6 : dato = 32'b01100110011001100110011001100110;
			11'h1c7 : dato = 32'b01100110011010001010001111110101;
			11'h1c8 : dato = 32'b11111111111111111111111111111111;
			11'h1c9 : dato = 32'b11111111111111111111111111111111;
			11'h1ca : dato = 32'b11111111111111111111111111111111;
			11'h1cb : dato = 32'b11111111111111111111111111111111;
			11'h1cc : dato = 32'b11111111111111111111111111111111;
			11'h1cd : dato = 32'b11111111111111111111111111111111;
			11'h1ce : dato = 32'b11111111111111111111111111111111;
			11'h1cf : dato = 32'b11111111111111111111111111111111;
			11'h1d0 : dato = 32'b11111111110001100110110101100110;
			11'h1d1 : dato = 32'b01100110011001100110011001100110;
			11'h1d2 : dato = 32'b01100110011001100110011001100110;
			11'h1d3 : dato = 32'b01100110011001100110011001100110;
			11'h1d4 : dato = 32'b01100110011001100110011001100110;
			11'h1d5 : dato = 32'b01100110011001100111010010011101;
			11'h1d6 : dato = 32'b10011000011011110110011001100110;
			11'h1d7 : dato = 32'b01100110011001100110011001100110;
			11'h1d8 : dato = 32'b01100110011001100110011001100110;
			11'h1d9 : dato = 32'b01100110011001100110011001100110;
			11'h1da : dato = 32'b01100110011001100110011001100110;
			11'h1db : dato = 32'b01100110011001100110011001110111;
			11'h1dc : dato = 32'b11010010111111111111111111111111;
			11'h1dd : dato = 32'b11111111111111111111111111111111;
			11'h1de : dato = 32'b11111111111111111111111111111111;
			11'h1df : dato = 32'b11111111111111111111111111111111;
			11'h1e0 : dato = 32'b11111111111111111111111111111111;
			11'h1e1 : dato = 32'b11111111111111111111111111111111;
			11'h1e2 : dato = 32'b11111111111111111111111111111111;
			11'h1e3 : dato = 32'b11111111111111111111111111111111;
			11'h1e4 : dato = 32'b11000001011001100110011001100110;
			11'h1e5 : dato = 32'b01100110011001100110011001100110;
			11'h1e6 : dato = 32'b01100110011001100110011001100110;
			11'h1e7 : dato = 32'b01100110011001100110011001100110;
			11'h1e8 : dato = 32'b01100110011001100110011001100110;
			11'h1e9 : dato = 32'b01100110011001100110011001100110;
			11'h1ea : dato = 32'b01100110011001100110011001100110;
			11'h1eb : dato = 32'b01100110011001100110011001100110;
			11'h1ec : dato = 32'b01100110011001100110011001100110;
			11'h1ed : dato = 32'b01100110011001100110011001100110;
			11'h1ee : dato = 32'b01100110011001100110011001100110;
			11'h1ef : dato = 32'b01100110011001100110011001100110;
			11'h1f0 : dato = 32'b01100110110000111111111111111111;
			11'h1f1 : dato = 32'b11111111111111111111111111111111;
			11'h1f2 : dato = 32'b11111111111111111111111111111111;
			11'h1f3 : dato = 32'b11111111111111111111111111111111;
			11'h1f4 : dato = 32'b11111111111111111111111111111111;
			11'h1f5 : dato = 32'b11111111111111111111111111111111;
			11'h1f6 : dato = 32'b11111111111111111111111111111111;
			11'h1f7 : dato = 32'b11111111111111111111111110111001;
			11'h1f8 : dato = 32'b01101000011001100110011001100110;
			11'h1f9 : dato = 32'b01100110011001100110011001100110;
			11'h1fa : dato = 32'b01100110011001100110011001100110;
			11'h1fb : dato = 32'b01100110011001100110011001100110;
			11'h1fc : dato = 32'b01100110011001100110011001100110;
			11'h1fd : dato = 32'b01100110011001100110011001100110;
			11'h1fe : dato = 32'b01100110011001100110011001100110;
			11'h1ff : dato = 32'b01100110011001100110011001100110;
			11'h200 : dato = 32'b01100110011001100110011001100110;
			11'h201 : dato = 32'b01100110011001100110011001100110;
			11'h202 : dato = 32'b01100110011001100110011001100110;
			11'h203 : dato = 32'b01100110011001100110011001100110;
			11'h204 : dato = 32'b01100110011010101101010011111111;
			11'h205 : dato = 32'b11111111111111111111111111111111;
			11'h206 : dato = 32'b11111111111111111111111111111111;
			11'h207 : dato = 32'b11111111111111111111111111111111;
			11'h208 : dato = 32'b11111111111111111111111111111111;
			11'h209 : dato = 32'b11111111111111111111111111111111;
			11'h20a : dato = 32'b11111111111111111111111111111111;
			11'h20b : dato = 32'b11111111111111111011011001100110;
			11'h20c : dato = 32'b01100110011001100110011001100110;
			11'h20d : dato = 32'b01100110011001100110011001100110;
			11'h20e : dato = 32'b01100110011001100110011001100110;
			11'h20f : dato = 32'b01100110011001100110011001100110;
			11'h210 : dato = 32'b01100110011001100110011001100110;
			11'h211 : dato = 32'b01100110011001100110011001100110;
			11'h212 : dato = 32'b01100110011001100110011001100110;
			11'h213 : dato = 32'b01100110011001100110011001100110;
			11'h214 : dato = 32'b01100110011001100110011001100110;
			11'h215 : dato = 32'b01100110011001100110011001100110;
			11'h216 : dato = 32'b01100110011001100110011001100110;
			11'h217 : dato = 32'b01100110011001100110011001100110;
			11'h218 : dato = 32'b01100110011001100110110111100110;
			11'h219 : dato = 32'b11111111111111111111111111111111;
			11'h21a : dato = 32'b11111111111111111111111111111111;
			11'h21b : dato = 32'b11111111111111111111111111111111;
			11'h21c : dato = 32'b11111111111111111111111111111111;
			11'h21d : dato = 32'b11111111111111111111111111111111;
			11'h21e : dato = 32'b11111111111111111111111111111111;
			11'h21f : dato = 32'b11111111110101000110011101100110;
			11'h220 : dato = 32'b01100110011001100110011001100110;
			11'h221 : dato = 32'b01100110011001100110011001100110;
			11'h222 : dato = 32'b01100110011001100110011001100110;
			11'h223 : dato = 32'b01100110011001100110011001100110;
			11'h224 : dato = 32'b01100110011001100110011001100110;
			11'h225 : dato = 32'b01100110011001100110011001100110;
			11'h226 : dato = 32'b01100110011001100110011001100110;
			11'h227 : dato = 32'b01100110011001100110011001100110;
			11'h228 : dato = 32'b01100110011001100110011001100110;
			11'h229 : dato = 32'b01100110011001100110011001100110;
			11'h22a : dato = 32'b01100110011001100110011001100110;
			11'h22b : dato = 32'b01100110011001100110011001100110;
			11'h22c : dato = 32'b01100110011001100110011010100010;
			11'h22d : dato = 32'b11111111111111111111111111111111;
			11'h22e : dato = 32'b11111111111111111111111111111111;
			11'h22f : dato = 32'b11111111111111111111111111111111;
			11'h230 : dato = 32'b11111111111111111111111111111111;
			11'h231 : dato = 32'b11111111111111111111111111111111;
			11'h232 : dato = 32'b11111111111111111111111111111111;
			11'h233 : dato = 32'b11111100011110000110011001100110;
			11'h234 : dato = 32'b01100110011001100110011001100110;
			11'h235 : dato = 32'b01100110011001100110011001100110;
			11'h236 : dato = 32'b01100110011001100110011001100110;
			11'h237 : dato = 32'b01100110011001100110011001100110;
			11'h238 : dato = 32'b01100110011001100110011001100110;
			11'h239 : dato = 32'b01100110011001100110011001100110;
			11'h23a : dato = 32'b01100110011001100110011001100110;
			11'h23b : dato = 32'b01100110011001100110011001100110;
			11'h23c : dato = 32'b01100110011001100110011001100110;
			11'h23d : dato = 32'b01100110011001100110011001100110;
			11'h23e : dato = 32'b01100110011001100110011001100110;
			11'h23f : dato = 32'b01100110011001100110011001100110;
			11'h240 : dato = 32'b01100110011001101010011111111110;
			11'h241 : dato = 32'b11111111111111111111111111111111;
			11'h242 : dato = 32'b11111111111111111111111111111111;
			11'h243 : dato = 32'b11111111111111111111111111111111;
			11'h244 : dato = 32'b11111111111111111111111111111111;
			11'h245 : dato = 32'b11111111111111111111111111111111;
			11'h246 : dato = 32'b11111111111111111111111111111111;
			11'h247 : dato = 32'b10111001011001100110011001100110;
			11'h248 : dato = 32'b01100110011001100110011001100110;
			11'h249 : dato = 32'b01100110011001100110011001100110;
			11'h24a : dato = 32'b01100110011001100110011001100110;
			11'h24b : dato = 32'b01100110011001100110011001100110;
			11'h24c : dato = 32'b01100110011001100110011001100110;
			11'h24d : dato = 32'b01100110011001100110011001100110;
			11'h24e : dato = 32'b01100110011001100110011001100110;
			11'h24f : dato = 32'b01100110011001100110011001100110;
			11'h250 : dato = 32'b01100110011001100110011001100110;
			11'h251 : dato = 32'b01100110011001100110011001100110;
			11'h252 : dato = 32'b01100110011001100110011001100110;
			11'h253 : dato = 32'b01100110011001100110011001100110;
			11'h254 : dato = 32'b01100111101110111111111111111111;
			11'h255 : dato = 32'b11111111111111111111111111111111;
			11'h256 : dato = 32'b11111111111111111111111111111111;
			11'h257 : dato = 32'b11111111111111111111111111111111;
			11'h258 : dato = 32'b11111111111111111111111111111111;
			11'h259 : dato = 32'b11111111111111111111111111111111;
			11'h25a : dato = 32'b11111111111111111111111111110000;
			11'h25b : dato = 32'b01101111011001100110011001100110;
			11'h25c : dato = 32'b01100110011001100110011001100110;
			11'h25d : dato = 32'b01100110011001100110011001100110;
			11'h25e : dato = 32'b01100110011001100110011001100110;
			11'h25f : dato = 32'b01100110011001100110011001100110;
			11'h260 : dato = 32'b01100110011001100110011001100110;
			11'h261 : dato = 32'b01100110011001100110011001100110;
			11'h262 : dato = 32'b01100110011001100110011001100110;
			11'h263 : dato = 32'b01100110011001100110011001100110;
			11'h264 : dato = 32'b01100110011001100110011001100110;
			11'h265 : dato = 32'b01100110011001100110011001100110;
			11'h266 : dato = 32'b01100110011001100110011001100110;
			11'h267 : dato = 32'b01100110011001100110011001110010;
			11'h268 : dato = 32'b11011101111111111111111111111111;
			11'h269 : dato = 32'b11111111111111111111111111111111;
			11'h26a : dato = 32'b11111111111111111111111111111111;
			11'h26b : dato = 32'b11111111111111111111111111111111;
			11'h26c : dato = 32'b11111111111111111111111111111111;
			11'h26d : dato = 32'b11111111111111111111111111111111;
			11'h26e : dato = 32'b11111111111111111111111110011000;
			11'h26f : dato = 32'b01100110011001100110011001100110;
			11'h270 : dato = 32'b01100110011001100110011001100110;
			11'h271 : dato = 32'b01100110011001100110011001100110;
			11'h272 : dato = 32'b01100110011001100110011001100110;
			11'h273 : dato = 32'b01100110011001100110011001100110;
			11'h274 : dato = 32'b01100110011001100110011001100110;
			11'h275 : dato = 32'b01100110011001100110011001100110;
			11'h276 : dato = 32'b01100110011001100110011001100110;
			11'h277 : dato = 32'b01100110011001100110011001100110;
			11'h278 : dato = 32'b01100110011001100110011001100110;
			11'h279 : dato = 32'b01100110011001100110011001100110;
			11'h27a : dato = 32'b01100110011001100110011001100110;
			11'h27b : dato = 32'b01100110011001100110101011011100;
			11'h27c : dato = 32'b11111111111111111111111111111111;
			11'h27d : dato = 32'b11111111111111111111111111111111;
			11'h27e : dato = 32'b11111111111111111111111111111111;
			11'h27f : dato = 32'b11111111111111111111111111111111;
			11'h280 : dato = 32'b11111111111111111111111111111111;
			11'h281 : dato = 32'b11111111111111111111111111111111;
			11'h282 : dato = 32'b11111111111111111110010001100110;
			11'h283 : dato = 32'b01100110011001100110011001100110;
			11'h284 : dato = 32'b01100110011001100110011001100110;
			11'h285 : dato = 32'b01100110011001100110011001100110;
			11'h286 : dato = 32'b01100110011001100110011001100110;
			11'h287 : dato = 32'b01100110011001100110011001100110;
			11'h288 : dato = 32'b01100110011001100110011001100110;
			11'h289 : dato = 32'b01100110011001100110011001100110;
			11'h28a : dato = 32'b01100110011001100110011001100110;
			11'h28b : dato = 32'b01100110011001100110011001100110;
			11'h28c : dato = 32'b01100110011001100110011001100110;
			11'h28d : dato = 32'b01100110011001100110011001100110;
			11'h28e : dato = 32'b01100110011001100110011001100110;
			11'h28f : dato = 32'b01100110011001101011100011111111;
			11'h290 : dato = 32'b11111111111111111111111111111111;
			11'h291 : dato = 32'b11111111111111111111111111111111;
			11'h292 : dato = 32'b11111111111111111111111111111111;
			11'h293 : dato = 32'b11111111111111111111111111111111;
			11'h294 : dato = 32'b11111111111111111111111111111111;
			11'h295 : dato = 32'b11111111111111111111111111111111;
			11'h296 : dato = 32'b11111111111111111011001001100110;
			11'h297 : dato = 32'b01100110011001100110011001100110;
			11'h298 : dato = 32'b01100110011001100110011001100110;
			11'h299 : dato = 32'b01100110011001100110011001100110;
			11'h29a : dato = 32'b01100110011001100110011001100110;
			11'h29b : dato = 32'b01100110011001100110011001100110;
			11'h29c : dato = 32'b01100110011001100110011001100110;
			11'h29d : dato = 32'b01100110011001100110011001100110;
			11'h29e : dato = 32'b01100110011001100110011001100110;
			11'h29f : dato = 32'b01100110011001100110011001100110;
			11'h2a0 : dato = 32'b01100110011001100110011001100110;
			11'h2a1 : dato = 32'b01100110011001100110011001100110;
			11'h2a2 : dato = 32'b01100110011001100110011001100110;
			11'h2a3 : dato = 32'b01100110011101011111110011111111;
			11'h2a4 : dato = 32'b11111111111111111111111111111111;
			11'h2a5 : dato = 32'b11111111111111111111111111111111;
			11'h2a6 : dato = 32'b11111111111111111111111111111111;
			11'h2a7 : dato = 32'b11111111111111111111111111111111;
			11'h2a8 : dato = 32'b11111111111111111111111111111111;
			11'h2a9 : dato = 32'b11111111111111111111111111111111;
			11'h2aa : dato = 32'b11111111111111111000011101100110;
			11'h2ab : dato = 32'b01100110011001100110011001100110;
			11'h2ac : dato = 32'b01100110011001100110011001100110;
			11'h2ad : dato = 32'b01100110011001100110011001100110;
			11'h2ae : dato = 32'b01100110011001100110011001100110;
			11'h2af : dato = 32'b01100110011001100110011001100110;
			11'h2b0 : dato = 32'b01100110011001100110011001100110;
			11'h2b1 : dato = 32'b01100110011001100110011001100110;
			11'h2b2 : dato = 32'b01100110011001100110011001100110;
			11'h2b3 : dato = 32'b01100110011001100110011001100110;
			11'h2b4 : dato = 32'b01100110011001100110011001100110;
			11'h2b5 : dato = 32'b01100110011001100110011001100110;
			11'h2b6 : dato = 32'b01100110011001100110011001100110;
			11'h2b7 : dato = 32'b01100110101110011111111111111111;
			11'h2b8 : dato = 32'b11111111111111111111111111111111;
			11'h2b9 : dato = 32'b11111111111111111111111111111111;
			11'h2ba : dato = 32'b11111111111111111111111111111111;
			11'h2bb : dato = 32'b11111111111111111111111111111111;
			11'h2bc : dato = 32'b11111111111111111111111111111111;
			11'h2bd : dato = 32'b11111111111111111111111111111111;
			11'h2be : dato = 32'b11111111111101000110011101100110;
			11'h2bf : dato = 32'b01100110011001100110011001100110;
			11'h2c0 : dato = 32'b01100110011001100110011001100110;
			11'h2c1 : dato = 32'b01100110011001100110011001100110;
			11'h2c2 : dato = 32'b01100110011001100110011001100110;
			11'h2c3 : dato = 32'b01100110011001100110011001100110;
			11'h2c4 : dato = 32'b01100110011001100110011001100110;
			11'h2c5 : dato = 32'b01100110011001100110011001100110;
			11'h2c6 : dato = 32'b01100110011001100110011001100110;
			11'h2c7 : dato = 32'b01100110011001100110011001100110;
			11'h2c8 : dato = 32'b01100110011001100110011001100110;
			11'h2c9 : dato = 32'b01100110011001100110011001100110;
			11'h2ca : dato = 32'b01100110011001100110011001100110;
			11'h2cb : dato = 32'b01101011111101011111111111111111;
			11'h2cc : dato = 32'b11111111111111111111111111111111;
			11'h2cd : dato = 32'b11111111111111111111111111111111;
			11'h2ce : dato = 32'b11111111111111111111111111111111;
			11'h2cf : dato = 32'b11111111111111111111111111111111;
			11'h2d0 : dato = 32'b11111111111111111111111111111111;
			11'h2d1 : dato = 32'b11111111111111111111111111111111;
			11'h2d2 : dato = 32'b11111111110100110110011001100110;
			11'h2d3 : dato = 32'b01100110011001100110011001100110;
			11'h2d4 : dato = 32'b01100110011001100110011001100110;
			11'h2d5 : dato = 32'b01100110011001100110011001100110;
			11'h2d6 : dato = 32'b01100110011001100110011001100110;
			11'h2d7 : dato = 32'b01100110011001100110011001100110;
			11'h2d8 : dato = 32'b01100110011001100110011001100110;
			11'h2d9 : dato = 32'b01100110011001100110011001100110;
			11'h2da : dato = 32'b01100110011001100110011001100110;
			11'h2db : dato = 32'b01100110011001100110011001100110;
			11'h2dc : dato = 32'b01100110011001100110011001100110;
			11'h2dd : dato = 32'b01100110011001100110011001100110;
			11'h2de : dato = 32'b01100110011001100110011001100110;
			11'h2df : dato = 32'b10010101111111111111111111111111;
			11'h2e0 : dato = 32'b11111111111111111111111111111111;
			11'h2e1 : dato = 32'b11111111111111111111111111111111;
			11'h2e2 : dato = 32'b11111111111111111111111111111111;
			11'h2e3 : dato = 32'b11111111111111111111111111111111;
			11'h2e4 : dato = 32'b11111111111111111111111111111111;
			11'h2e5 : dato = 32'b11111111111111111111111111111111;
			11'h2e6 : dato = 32'b11111111101110010110011001100110;
			11'h2e7 : dato = 32'b01100110011001100110011001100110;
			11'h2e8 : dato = 32'b01100110011001100110011001100110;
			11'h2e9 : dato = 32'b01100110011001100110011001100110;
			11'h2ea : dato = 32'b01100110011001100110011001100110;
			11'h2eb : dato = 32'b01100110011001100110011001100110;
			11'h2ec : dato = 32'b01100110011001100110011001100110;
			11'h2ed : dato = 32'b01100110011001100110011001100110;
			11'h2ee : dato = 32'b01100110011001100110011001100110;
			11'h2ef : dato = 32'b01100110011001100110011001100110;
			11'h2f0 : dato = 32'b01100110011001100110011001100110;
			11'h2f1 : dato = 32'b01100110011001100110011001100110;
			11'h2f2 : dato = 32'b01100110011001100110011001100110;
			11'h2f3 : dato = 32'b10111000111111111111111111111111;
			11'h2f4 : dato = 32'b11111111111111111111111111111111;
			11'h2f5 : dato = 32'b11111111111111111111111111111111;
			11'h2f6 : dato = 32'b11111111111111111111111111111111;
			11'h2f7 : dato = 32'b11111111111111111111111111111111;
			11'h2f8 : dato = 32'b11111111111111111111111111111111;
			11'h2f9 : dato = 32'b11111111111111111111111111111111;
			11'h2fa : dato = 32'b11111111101001110110011001100110;
			11'h2fb : dato = 32'b01100110011001100110011001100110;
			11'h2fc : dato = 32'b01100110011001100110011001100110;
			11'h2fd : dato = 32'b01100110011001100110011001100110;
			11'h2fe : dato = 32'b01100110011001100110011001100110;
			11'h2ff : dato = 32'b01100110011001100110011001100110;
			11'h300 : dato = 32'b01100110011001100110011001100110;
			11'h301 : dato = 32'b01100110011001100110011001100110;
			11'h302 : dato = 32'b01100110011001100110011001100110;
			11'h303 : dato = 32'b01100110011001100110011001100110;
			11'h304 : dato = 32'b01100110011001100110011001100110;
			11'h305 : dato = 32'b01100110011001100110011001100110;
			11'h306 : dato = 32'b01100110011001100110011001100110;
			11'h307 : dato = 32'b11010010111111111111111111111111;
			11'h308 : dato = 32'b11111111111111111111111111111111;
			11'h309 : dato = 32'b11111111111111111111111111111111;
			11'h30a : dato = 32'b11111111111111111111111111111111;
			11'h30b : dato = 32'b11111111111111111111111111111111;
			11'h30c : dato = 32'b11111111111111111111111111111111;
			11'h30d : dato = 32'b11111111111111111111111111111111;
			11'h30e : dato = 32'b11111111100100110110011001100110;
			11'h30f : dato = 32'b01100110011001100110011001100110;
			11'h310 : dato = 32'b01100110011001100110011001100110;
			11'h311 : dato = 32'b01100110011001100110011001100110;
			11'h312 : dato = 32'b01100110011001100110011001100110;
			11'h313 : dato = 32'b01100110011001100110011001100110;
			11'h314 : dato = 32'b01100110011001100110011001100110;
			11'h315 : dato = 32'b01100110011001100110011001100110;
			11'h316 : dato = 32'b01100110011001100110011001100110;
			11'h317 : dato = 32'b01100110011001100110011001100110;
			11'h318 : dato = 32'b01100110011001100110011001100110;
			11'h319 : dato = 32'b01100110011001100110011001100110;
			11'h31a : dato = 32'b01100110011001100110011001100110;
			11'h31b : dato = 32'b11101010111111111111111111111111;
			11'h31c : dato = 32'b11111111111111111111111111111111;
			11'h31d : dato = 32'b11111111111111111111111111111111;
			11'h31e : dato = 32'b11111111111111111111111111111111;
			11'h31f : dato = 32'b11111111111111111111111111111111;
			11'h320 : dato = 32'b11111111111111111111111111111111;
			11'h321 : dato = 32'b11111111111111111111111111111111;
			11'h322 : dato = 32'b11111111100001110110011001100110;
			11'h323 : dato = 32'b01100110011001100110011001100110;
			11'h324 : dato = 32'b01100110011001100110011001100110;
			11'h325 : dato = 32'b01100110011001100110011001100110;
			11'h326 : dato = 32'b01100110011001100110011001100110;
			11'h327 : dato = 32'b01100110011001100110011001100110;
			11'h328 : dato = 32'b01100110011001100110011001100110;
			11'h329 : dato = 32'b01100110011001100110011001100110;
			11'h32a : dato = 32'b01100110011001100110011001100110;
			11'h32b : dato = 32'b01100110011001100110011001100110;
			11'h32c : dato = 32'b01100110011001100110011001100110;
			11'h32d : dato = 32'b01100110011001100110011001100110;
			11'h32e : dato = 32'b01100110011001100110011001100110;
			11'h32f : dato = 32'b11110111111111111111111111111111;
			11'h330 : dato = 32'b11111111111111111111111111111111;
			11'h331 : dato = 32'b11111111111111111111111111111111;
			11'h332 : dato = 32'b11111111111111111111111111111111;
			11'h333 : dato = 32'b11111111111111111111111111111111;
			11'h334 : dato = 32'b11111111111111111111111111111111;
			11'h335 : dato = 32'b11111111111111111111111111111111;
			11'h336 : dato = 32'b11111111100001000110011001100110;
			11'h337 : dato = 32'b01100110011001100110011001100110;
			11'h338 : dato = 32'b01100110011001100110011001100110;
			11'h339 : dato = 32'b01100110011001100110011001100110;
			11'h33a : dato = 32'b01100110011001100110011001100110;
			11'h33b : dato = 32'b01100110011001100110011001100110;
			11'h33c : dato = 32'b01100110011001100110011001100110;
			11'h33d : dato = 32'b01100110011001100110011001100110;
			11'h33e : dato = 32'b01100110011001100110011001100110;
			11'h33f : dato = 32'b01100110011001100110011001100110;
			11'h340 : dato = 32'b01100110011001100110011001100110;
			11'h341 : dato = 32'b01100110011001100110011001100110;
			11'h342 : dato = 32'b01100110011001100110011001100110;
			11'h343 : dato = 32'b11111000111111111111111111111111;
			11'h344 : dato = 32'b11111111111111111111111111111111;
			11'h345 : dato = 32'b11111111111111111111111111111111;
			11'h346 : dato = 32'b11111111111111111111111111111111;
			11'h347 : dato = 32'b11111111111111111111111111111111;
			11'h348 : dato = 32'b11111111111111111111111111111111;
			11'h349 : dato = 32'b11111111111111111111111111111111;
			11'h34a : dato = 32'b11111111100000110110011001100110;
			11'h34b : dato = 32'b01100110011001100110011001100110;
			11'h34c : dato = 32'b01100110011001100110011001100110;
			11'h34d : dato = 32'b01100110011001100110011001100110;
			11'h34e : dato = 32'b01100110011001100110011001100110;
			11'h34f : dato = 32'b01100110011001100110011001100110;
			11'h350 : dato = 32'b01100110011001100110011001100110;
			11'h351 : dato = 32'b01100110011001100110011001100110;
			11'h352 : dato = 32'b01100110011001100110011001100110;
			11'h353 : dato = 32'b01100110011001100110011001100110;
			11'h354 : dato = 32'b01100110011001100110011001100110;
			11'h355 : dato = 32'b01100110011001100110011001100110;
			11'h356 : dato = 32'b01100110011001100110011001100110;
			11'h357 : dato = 32'b11110111111111111111111111111111;
			11'h358 : dato = 32'b11111111111111111111111111111111;
			11'h359 : dato = 32'b11111111111111111111111111111111;
			11'h35a : dato = 32'b11111111111111111111111111111111;
			11'h35b : dato = 32'b11111111111111111111111111111111;
			11'h35c : dato = 32'b11111111111111111111111111111111;
			11'h35d : dato = 32'b11111111111111111111111111111111;
			11'h35e : dato = 32'b11111111100001000110011001100110;
			11'h35f : dato = 32'b01100110011001100110011001100110;
			11'h360 : dato = 32'b01100110011001100110011001100110;
			11'h361 : dato = 32'b01100110011001100110011001100110;
			11'h362 : dato = 32'b01100110011001100110011001100110;
			11'h363 : dato = 32'b01100110011001100110011001100110;
			11'h364 : dato = 32'b01100110011001100110011001100110;
			11'h365 : dato = 32'b01100110011001100110011001100110;
			11'h366 : dato = 32'b01100110011001100110011001100110;
			11'h367 : dato = 32'b01100110011001100110011001100110;
			11'h368 : dato = 32'b01100110011001100110011001100110;
			11'h369 : dato = 32'b01100110011001100110011001100110;
			11'h36a : dato = 32'b01100110011001100110011001100110;
			11'h36b : dato = 32'b11110000111111111111111111111111;
			11'h36c : dato = 32'b11111111111111111111111111111111;
			11'h36d : dato = 32'b11111111111111111111111111111111;
			11'h36e : dato = 32'b11111111111111111111111111111111;
			11'h36f : dato = 32'b11111111111111111111111111111111;
			11'h370 : dato = 32'b11111111111111111111111111111111;
			11'h371 : dato = 32'b11111111111111111111111111111111;
			11'h372 : dato = 32'b11111111100001100110011001100110;
			11'h373 : dato = 32'b01100110011001100110011001100110;
			11'h374 : dato = 32'b01100110011001100110011001100110;
			11'h375 : dato = 32'b01100110011001100110011001100110;
			11'h376 : dato = 32'b01100110011001100110011001100110;
			11'h377 : dato = 32'b01100110011001100110011001100110;
			11'h378 : dato = 32'b01100110011001100110011001100110;
			11'h379 : dato = 32'b01100110011001100110011001100110;
			11'h37a : dato = 32'b01100110011001100110011001100110;
			11'h37b : dato = 32'b01100110011001100110011001100110;
			11'h37c : dato = 32'b01100110011001100110011001100110;
			11'h37d : dato = 32'b01100110011001100110011001100110;
			11'h37e : dato = 32'b01100110011001100110011001100110;
			11'h37f : dato = 32'b11011010111111111111111111111111;
			11'h380 : dato = 32'b11111111111111111111111111111111;
			11'h381 : dato = 32'b11111111111111111111111111111111;
			11'h382 : dato = 32'b11111111111111111111111111111111;
			11'h383 : dato = 32'b11111111111111111111111111111111;
			11'h384 : dato = 32'b11111111111111111111111111111111;
			11'h385 : dato = 32'b11111111111111111111111111111111;
			11'h386 : dato = 32'b11111111100100000110011001100110;
			11'h387 : dato = 32'b01100110011001100110011001100110;
			11'h388 : dato = 32'b01100110011001100110011001100110;
			11'h389 : dato = 32'b01100110011001100110011001100110;
			11'h38a : dato = 32'b01100110011001100110011001100110;
			11'h38b : dato = 32'b01100110011001100110011001100110;
			11'h38c : dato = 32'b01100110011001100110011001100110;
			11'h38d : dato = 32'b01100110011001100110011001100110;
			11'h38e : dato = 32'b01100110011001100110011001100110;
			11'h38f : dato = 32'b01100110011001100110011001100110;
			11'h390 : dato = 32'b01100110011001100110011001100110;
			11'h391 : dato = 32'b01100110011001100110011001100110;
			11'h392 : dato = 32'b01100110011001100110011001100110;
			11'h393 : dato = 32'b10111101111111111111111111111111;
			11'h394 : dato = 32'b11111111111111111111111111111111;
			11'h395 : dato = 32'b11111111111111111111111111111111;
			11'h396 : dato = 32'b11111111111111111111111111111111;
			11'h397 : dato = 32'b11111111111111111111111111111111;
			11'h398 : dato = 32'b11111111111111111111111111111111;
			11'h399 : dato = 32'b11111111111111111111111111111111;
			11'h39a : dato = 32'b11111111100111010110011001100110;
			11'h39b : dato = 32'b01100110011001100110011001100110;
			11'h39c : dato = 32'b01100110011001100110011001100110;
			11'h39d : dato = 32'b01100110011001100110011001100110;
			11'h39e : dato = 32'b01100110011001100110011001100110;
			11'h39f : dato = 32'b01100110011001100110011001100110;
			11'h3a0 : dato = 32'b01100110011001100110011001100110;
			11'h3a1 : dato = 32'b01100110011001100110011001100110;
			11'h3a2 : dato = 32'b01100110011001100110011001100110;
			11'h3a3 : dato = 32'b01100110011001100110011001100110;
			11'h3a4 : dato = 32'b01100110011001100110011001100110;
			11'h3a5 : dato = 32'b01100110011001100110011001100110;
			11'h3a6 : dato = 32'b01100110011001100110011001100110;
			11'h3a7 : dato = 32'b10011000111111111111111111111111;
			11'h3a8 : dato = 32'b11111111111111111111111111111111;
			11'h3a9 : dato = 32'b11111111111111111111111111111111;
			11'h3aa : dato = 32'b11111111111111111111111111111111;
			11'h3ab : dato = 32'b11111111111111111111111111111111;
			11'h3ac : dato = 32'b11111111111111111111111111111111;
			11'h3ad : dato = 32'b11111111111111111111111111111111;
			11'h3ae : dato = 32'b11111111101011000110011001100110;
			11'h3af : dato = 32'b01100110011001100110011001100110;
			11'h3b0 : dato = 32'b01100110011001100110011001100110;
			11'h3b1 : dato = 32'b01100110011001100110011001100110;
			11'h3b2 : dato = 32'b01100110011001100110011001100110;
			11'h3b3 : dato = 32'b01100110011001100110011001100110;
			11'h3b4 : dato = 32'b01100110011001100110011001100110;
			11'h3b5 : dato = 32'b01100110011001100110011001100110;
			11'h3b6 : dato = 32'b01100110011001100110011001100110;
			11'h3b7 : dato = 32'b01100110011001100110011001100110;
			11'h3b8 : dato = 32'b01100110011001100110011001100110;
			11'h3b9 : dato = 32'b01100110011001100110011001100110;
			11'h3ba : dato = 32'b01100110011001100110011001100110;
			11'h3bb : dato = 32'b01110000111110101111111111111111;
			11'h3bc : dato = 32'b11111111111111111111111111111111;
			11'h3bd : dato = 32'b11111111111111111111111111111111;
			11'h3be : dato = 32'b11111111111111111111111111111111;
			11'h3bf : dato = 32'b11111111111111111111111111111111;
			11'h3c0 : dato = 32'b11111111111111111111111111111111;
			11'h3c1 : dato = 32'b11111111111111111111111111111111;
			11'h3c2 : dato = 32'b11111111110000010110011001100110;
			11'h3c3 : dato = 32'b01100110011001100110011001100110;
			11'h3c4 : dato = 32'b01100110011001100110011001100110;
			11'h3c5 : dato = 32'b01100110011001100110011001100110;
			11'h3c6 : dato = 32'b01100110011001100110011001100110;
			11'h3c7 : dato = 32'b01100110011001100110011001100110;
			11'h3c8 : dato = 32'b01100110011001100110011001100110;
			11'h3c9 : dato = 32'b01100110011001100110011001100110;
			11'h3ca : dato = 32'b01100110011001100110011001100110;
			11'h3cb : dato = 32'b01100110011001100110011001100110;
			11'h3cc : dato = 32'b01100110011001100110011001100110;
			11'h3cd : dato = 32'b01100110011001100110011001100110;
			11'h3ce : dato = 32'b01100110011001100110011001100110;
			11'h3cf : dato = 32'b01100110110001011111111111111111;
			11'h3d0 : dato = 32'b11111111111111111111111111111111;
			11'h3d1 : dato = 32'b11111111111111111111111111111111;
			11'h3d2 : dato = 32'b11111111111111111111111111111111;
			11'h3d3 : dato = 32'b11111111111111111111111111111111;
			11'h3d4 : dato = 32'b11111111111111111111111111111111;
			11'h3d5 : dato = 32'b11111111111111111111111111111111;
			11'h3d6 : dato = 32'b11111111110110100110011001100110;
			11'h3d7 : dato = 32'b01100110011001100110011001100110;
			11'h3d8 : dato = 32'b01100110011001100110011001100110;
			11'h3d9 : dato = 32'b01100110011001100110011001100110;
			11'h3da : dato = 32'b01100110011001100110011001100110;
			11'h3db : dato = 32'b01100110011001100110011001100110;
			11'h3dc : dato = 32'b01100110011001100110011001100110;
			11'h3dd : dato = 32'b01100110011001100110011001100110;
			11'h3de : dato = 32'b01100110011001100110011001100110;
			11'h3df : dato = 32'b01100110011001100110011001100110;
			11'h3e0 : dato = 32'b01100110011001100110011001100110;
			11'h3e1 : dato = 32'b01100110011001100110011001100110;
			11'h3e2 : dato = 32'b01100110011001100110011001100110;
			11'h3e3 : dato = 32'b01100110011111001111110011111111;
			11'h3e4 : dato = 32'b11111111111111111111111111111111;
			11'h3e5 : dato = 32'b11111111111111111111111111111111;
			11'h3e6 : dato = 32'b11111111111111111111111111111111;
			11'h3e7 : dato = 32'b11111111111111111111111111111111;
			11'h3e8 : dato = 32'b11111111111111111111111111111111;
			11'h3e9 : dato = 32'b11111111111111111111111111111111;
			11'h3ea : dato = 32'b11111111111101100110011101100110;
			11'h3eb : dato = 32'b01100110011001100110011001100110;
			11'h3ec : dato = 32'b01100110011001100110011001100110;
			11'h3ed : dato = 32'b01100110011001100110011001100110;
			11'h3ee : dato = 32'b01100110011001100110011001100110;
			11'h3ef : dato = 32'b01100110011001100110011001100110;
			11'h3f0 : dato = 32'b01100110011001100110011001100110;
			11'h3f1 : dato = 32'b01100110011001100110011001100110;
			11'h3f2 : dato = 32'b01100110011001100110011001100110;
			11'h3f3 : dato = 32'b01100110011001100110011001100110;
			11'h3f4 : dato = 32'b01100110011001100110011001100110;
			11'h3f5 : dato = 32'b01100110011001100110011001100110;
			11'h3f6 : dato = 32'b01100110011001100110011001100110;
			11'h3f7 : dato = 32'b01100110011001101011011111111111;
			11'h3f8 : dato = 32'b11111111111111111111111111111111;
			11'h3f9 : dato = 32'b11111111111111111111111111111111;
			11'h3fa : dato = 32'b11111111111111111111111111111111;
			11'h3fb : dato = 32'b11111111111111111111111111111111;
			11'h3fc : dato = 32'b11111111111111111111111111111111;
			11'h3fd : dato = 32'b11111111111111111111111111111111;
			11'h3fe : dato = 32'b11111111111111110111101101100110;
			11'h3ff : dato = 32'b01100110011001100110011001100110;
			11'h400 : dato = 32'b01100110011001100110011001100110;
			11'h401 : dato = 32'b01100110011001100110011001100110;
			11'h402 : dato = 32'b01100110011001100110011001100110;
			11'h403 : dato = 32'b01100110011001100110011001100110;
			11'h404 : dato = 32'b01100110011001100110011001100110;
			11'h405 : dato = 32'b01100110011001100110011001100110;
			11'h406 : dato = 32'b01100110011001100110011001100110;
			11'h407 : dato = 32'b01100110011001100110011001100110;
			11'h408 : dato = 32'b01100110011001100110011001100110;
			11'h409 : dato = 32'b01100110011001100110011001100110;
			11'h40a : dato = 32'b01100110011001100110011001100110;
			11'h40b : dato = 32'b01100110011001100110110011101110;
			11'h40c : dato = 32'b11111111111111111111111111111111;
			11'h40d : dato = 32'b11111111111111111111111111111111;
			11'h40e : dato = 32'b11111111111111111111111111111111;
			11'h40f : dato = 32'b11111111111111111111111111111111;
			11'h410 : dato = 32'b11111111111111111111111111111111;
			11'h411 : dato = 32'b11111111111111111111111111111111;
			11'h412 : dato = 32'b11111111111111111001101001100110;
			11'h413 : dato = 32'b01100110011001100110011001100110;
			11'h414 : dato = 32'b01100110011001100110011001100110;
			11'h415 : dato = 32'b01100110011001100110011001100110;
			11'h416 : dato = 32'b01100110011001100110011001100110;
			11'h417 : dato = 32'b01100110011001100110011001100110;
			11'h418 : dato = 32'b01100110011001100110011001100110;
			11'h419 : dato = 32'b01100110011001100110011001100110;
			11'h41a : dato = 32'b01100110011001100110011001100110;
			11'h41b : dato = 32'b01100110011001100110011001100110;
			11'h41c : dato = 32'b01100110011001100110011001100110;
			11'h41d : dato = 32'b01100110011001100110011001100110;
			11'h41e : dato = 32'b01100110011001100110011001100110;
			11'h41f : dato = 32'b01100110011001100110011010001101;
			11'h420 : dato = 32'b11111010111111111111111111111111;
			11'h421 : dato = 32'b11111111111111111111111111111111;
			11'h422 : dato = 32'b11111111111111111111111111111111;
			11'h423 : dato = 32'b11111111111111111111111111111111;
			11'h424 : dato = 32'b11111111111111111111111111111111;
			11'h425 : dato = 32'b11111111111111111111111111111111;
			11'h426 : dato = 32'b11111111111111111100001001100110;
			11'h427 : dato = 32'b01100110011001100110011001100110;
			11'h428 : dato = 32'b01100110011001100110011001100110;
			11'h429 : dato = 32'b01100110011001100110011001100110;
			11'h42a : dato = 32'b01100110011001100110011001100110;
			11'h42b : dato = 32'b01100110011001100110011001100110;
			11'h42c : dato = 32'b01100110011001100110011001100110;
			11'h42d : dato = 32'b01100110011001100110011001100110;
			11'h42e : dato = 32'b01100110011001100110011001100110;
			11'h42f : dato = 32'b01100110011001100110011001100110;
			11'h430 : dato = 32'b01100110011001100110011001100110;
			11'h431 : dato = 32'b01100110011001100110011001100110;
			11'h432 : dato = 32'b01100110011001100110011001100110;
			11'h433 : dato = 32'b01100110011001100110011001100110;
			11'h434 : dato = 32'b10000100111011101111111111111111;
			11'h435 : dato = 32'b11111111111111111111111111111111;
			11'h436 : dato = 32'b11111111111111111111111111111111;
			11'h437 : dato = 32'b11111111111111111111111111111111;
			11'h438 : dato = 32'b11111111111111111111111111111111;
			11'h439 : dato = 32'b11111111111111111111111111111111;
			11'h43a : dato = 32'b11111111111111111110111001100110;
			11'h43b : dato = 32'b01100110011001100110011001100110;
			11'h43c : dato = 32'b01100110011001100110011001100110;
			11'h43d : dato = 32'b01100110011001100110011001100110;
			11'h43e : dato = 32'b01100110011001100110011001100110;
			11'h43f : dato = 32'b01100110011001100110011001100110;
			11'h440 : dato = 32'b01100110011001100110011001100110;
			11'h441 : dato = 32'b01100110011001100110011001100110;
			11'h442 : dato = 32'b01100110011001100110011001100110;
			11'h443 : dato = 32'b01100110011001100110011001100110;
			11'h444 : dato = 32'b01100110011001100110011001100110;
			11'h445 : dato = 32'b01100110011001100110011001100110;
			11'h446 : dato = 32'b01100110011001100110011001100110;
			11'h447 : dato = 32'b01100110011001100110011001100110;
			11'h448 : dato = 32'b01100110011101101101111011111111;
			11'h449 : dato = 32'b11111111111111111111111111111111;
			11'h44a : dato = 32'b11111111111111111111111111111111;
			11'h44b : dato = 32'b11111111111111111111111111111111;
			11'h44c : dato = 32'b11111111111111111111111111111111;
			11'h44d : dato = 32'b11111111111111111111111111111111;
			11'h44e : dato = 32'b11111111111111111111111110000101;
			11'h44f : dato = 32'b01100110011001100110011001100110;
			11'h450 : dato = 32'b01100110011001100110011001100110;
			11'h451 : dato = 32'b01100110011001100110011001100110;
			11'h452 : dato = 32'b01100110011001100110011001100110;
			11'h453 : dato = 32'b01100110011001100110011001100110;
			11'h454 : dato = 32'b01100110011001100110011001100110;
			11'h455 : dato = 32'b01100110011001100110011001100110;
			11'h456 : dato = 32'b01100110011001100110011001100110;
			11'h457 : dato = 32'b01100110011001100110011001100110;
			11'h458 : dato = 32'b01100110011001100110011001100110;
			11'h459 : dato = 32'b01100110011001100110011001100110;
			11'h45a : dato = 32'b01100110011001100110011001100110;
			11'h45b : dato = 32'b01100110011001100110011001100110;
			11'h45c : dato = 32'b01100110011001100110101011001001;
			11'h45d : dato = 32'b11111111111111111111111111111111;
			11'h45e : dato = 32'b11111111111111111111111111111111;
			11'h45f : dato = 32'b11111111111111111111111111111111;
			11'h460 : dato = 32'b11111111111111111111111111111111;
			11'h461 : dato = 32'b11111111111111111111111111111111;
			11'h462 : dato = 32'b11111111111111111111111111000000;
			11'h463 : dato = 32'b01100110011001100110011001100110;
			11'h464 : dato = 32'b01100110011001100110011001100110;
			11'h465 : dato = 32'b01100110011001100110011001100110;
			11'h466 : dato = 32'b01100110011001100110011001100110;
			11'h467 : dato = 32'b01100110011001100110011001100110;
			11'h468 : dato = 32'b01100110011001100110011001100110;
			11'h469 : dato = 32'b01100110011001100110011001100110;
			11'h46a : dato = 32'b01100110011001100110011001100110;
			11'h46b : dato = 32'b01100110011001100110011001100110;
			11'h46c : dato = 32'b01100110011001100110011001100110;
			11'h46d : dato = 32'b01100110011001100110011001100110;
			11'h46e : dato = 32'b01100110011001100110011001100110;
			11'h46f : dato = 32'b01100110011001100110011001100110;
			11'h470 : dato = 32'b01100110011001100110011001100110;
			11'h471 : dato = 32'b10001110110101011111111111111111;
			11'h472 : dato = 32'b11111111111111111111111111111111;
			11'h473 : dato = 32'b11111111111111111111111111111111;
			11'h474 : dato = 32'b11111111111111111111111111111111;
			11'h475 : dato = 32'b11111111111111111111111111111111;
			11'h476 : dato = 32'b11111111111111111111111111111010;
			11'h477 : dato = 32'b01110001011001100110011001100110;
			11'h478 : dato = 32'b01100110011001100110011001100110;
			11'h479 : dato = 32'b01100110011001100110011001100110;
			11'h47a : dato = 32'b01100110011001100110011001100110;
			11'h47b : dato = 32'b01100110011001100110011001100110;
			11'h47c : dato = 32'b01100110011001100110011001100110;
			11'h47d : dato = 32'b01100110011001100110011001100110;
			11'h47e : dato = 32'b01100110011001100110011001100110;
			11'h47f : dato = 32'b01100110011001100110011001100110;
			11'h480 : dato = 32'b01100110011001100110011001100110;
			11'h481 : dato = 32'b01100110011001100110011001100110;
			11'h482 : dato = 32'b01100110011001100110011001100110;
			11'h483 : dato = 32'b01100110011001100110011001100110;
			11'h484 : dato = 32'b01100110011001100110011001100110;
			11'h485 : dato = 32'b01100110100100001111111111111111;
			11'h486 : dato = 32'b11111111111111111111111111111111;
			11'h487 : dato = 32'b11111111111111111111111111111111;
			11'h488 : dato = 32'b11111111111111111111111111111111;
			11'h489 : dato = 32'b11111111111111111111111111111111;
			11'h48a : dato = 32'b11111111111111111111111111111111;
			11'h48b : dato = 32'b10100111011001100110011001100110;
			11'h48c : dato = 32'b01100110011001100110011001100110;
			11'h48d : dato = 32'b01100110011001100110011001100110;
			11'h48e : dato = 32'b01100110011001100110011001100110;
			11'h48f : dato = 32'b01100110011001100110011001100110;
			11'h490 : dato = 32'b01100110011001100110011001100110;
			11'h491 : dato = 32'b01100110011001100110011001100110;
			11'h492 : dato = 32'b01100110011001100110011001100110;
			11'h493 : dato = 32'b01100110011001100110011001100110;
			11'h494 : dato = 32'b01100110011001100110011001100110;
			11'h495 : dato = 32'b01100110011001100110011001100110;
			11'h496 : dato = 32'b01100110011001100110011001100110;
			11'h497 : dato = 32'b01100110011001100110011001100110;
			11'h498 : dato = 32'b01100110011001100110011001100110;
			11'h499 : dato = 32'b01100110110001001111111111111111;
			11'h49a : dato = 32'b11111111111111111111111111111111;
			11'h49b : dato = 32'b11111111111111111111111111111111;
			11'h49c : dato = 32'b11111111111111111111111111111111;
			11'h49d : dato = 32'b11111111111111111111111111111111;
			11'h49e : dato = 32'b11111111111111111111111111111111;
			11'h49f : dato = 32'b11011101011001100110011001100110;
			11'h4a0 : dato = 32'b01100110011001100110011001100110;
			11'h4a1 : dato = 32'b01100110011001100110011001100110;
			11'h4a2 : dato = 32'b01100110011001100110011001100110;
			11'h4a3 : dato = 32'b01100110011001100110011001100110;
			11'h4a4 : dato = 32'b01100110011001100110011001100110;
			11'h4a5 : dato = 32'b01100110011001100110011001100110;
			11'h4a6 : dato = 32'b01100110011001100110011001100110;
			11'h4a7 : dato = 32'b01100110011001100110011001100110;
			11'h4a8 : dato = 32'b01100110011001100110011001100110;
			11'h4a9 : dato = 32'b01100110011001100110011001100110;
			11'h4aa : dato = 32'b01100110011001100110011001100110;
			11'h4ab : dato = 32'b01100110011001100110011001100110;
			11'h4ac : dato = 32'b01100110011001100110011001100110;
			11'h4ad : dato = 32'b01101001111101011111111111111111;
			11'h4ae : dato = 32'b11111111111111111111111111111111;
			11'h4af : dato = 32'b11111111111111111111111111111111;
			11'h4b0 : dato = 32'b11111111111111111111111111111111;
			11'h4b1 : dato = 32'b11111111111111111111111111111111;
			11'h4b2 : dato = 32'b11111111111111111111111111111111;
			11'h4b3 : dato = 32'b11111110011111100110011001100110;
			11'h4b4 : dato = 32'b01100110011001100110011001100110;
			11'h4b5 : dato = 32'b01100110011001100110011001100110;
			11'h4b6 : dato = 32'b01100110011001100110011001100110;
			11'h4b7 : dato = 32'b01100110011001100110011001100110;
			11'h4b8 : dato = 32'b01100110011001100110011001100110;
			11'h4b9 : dato = 32'b01100110011001100110011001100110;
			11'h4ba : dato = 32'b01100110011001100110011001100110;
			11'h4bb : dato = 32'b01100110011001100110011001100110;
			11'h4bc : dato = 32'b01100110011001100110011001100110;
			11'h4bd : dato = 32'b01100110011001100110011001100110;
			11'h4be : dato = 32'b01100110011001100110011001100110;
			11'h4bf : dato = 32'b01100110011001100110011001100110;
			11'h4c0 : dato = 32'b01100110011001100110011001100110;
			11'h4c1 : dato = 32'b10100011111111111111111111111111;
			11'h4c2 : dato = 32'b11111111111111111111111111111111;
			11'h4c3 : dato = 32'b11111111111111111111111111111111;
			11'h4c4 : dato = 32'b11111111111111111111111111111111;
			11'h4c5 : dato = 32'b11111111111111111111111111111111;
			11'h4c6 : dato = 32'b11111111111111111111111111111111;
			11'h4c7 : dato = 32'b11111111110000110110011001100110;
			11'h4c8 : dato = 32'b01100110011001100110011001100110;
			11'h4c9 : dato = 32'b01100110011001100110011001100110;
			11'h4ca : dato = 32'b01100110011001100110011001100110;
			11'h4cb : dato = 32'b01100110011001100110011001100110;
			11'h4cc : dato = 32'b01100110011001100110011001100110;
			11'h4cd : dato = 32'b01100110011001100110011001100110;
			11'h4ce : dato = 32'b01100110011001100110011001100110;
			11'h4cf : dato = 32'b01100110011001100110011001100110;
			11'h4d0 : dato = 32'b01100110011001100110011001100110;
			11'h4d1 : dato = 32'b01100110011001100110011001100110;
			11'h4d2 : dato = 32'b01100110011001100110011001100110;
			11'h4d3 : dato = 32'b01100110011001100110011001100110;
			11'h4d4 : dato = 32'b01100110011001100110011001101110;
			11'h4d5 : dato = 32'b11110010111111111111111111111111;
			11'h4d6 : dato = 32'b11111111111111111111111111111111;
			11'h4d7 : dato = 32'b11111111111111111111111111111111;
			11'h4d8 : dato = 32'b11111111111111111111111111111111;
			11'h4d9 : dato = 32'b11111111111111111111111111111111;
			11'h4da : dato = 32'b11111111111111111111111111111111;
			11'h4db : dato = 32'b11111111111111000111100101100110;
			11'h4dc : dato = 32'b01100110011001100110011001100110;
			11'h4dd : dato = 32'b01100110011001100110011001100110;
			11'h4de : dato = 32'b01100110011001100110011001100110;
			11'h4df : dato = 32'b01100110011001100110011001100110;
			11'h4e0 : dato = 32'b01100110011001100110011001100110;
			11'h4e1 : dato = 32'b01100110011001100110011001100110;
			11'h4e2 : dato = 32'b01100110011001100110011001100110;
			11'h4e3 : dato = 32'b01100110011001100110011001100110;
			11'h4e4 : dato = 32'b01100110011001100110011001100110;
			11'h4e5 : dato = 32'b01100110011001100110011001100110;
			11'h4e6 : dato = 32'b01100110011001100110011001100110;
			11'h4e7 : dato = 32'b01100110011001100110011001100110;
			11'h4e8 : dato = 32'b01100110011001100110011010101011;
			11'h4e9 : dato = 32'b11111111111111111111111111111111;
			11'h4ea : dato = 32'b11111111111111111111111111111111;
			11'h4eb : dato = 32'b11111111111111111111111111111111;
			11'h4ec : dato = 32'b11111111111111111111111111111111;
			11'h4ed : dato = 32'b11111111111111111111111111111111;
			11'h4ee : dato = 32'b11111111111111111111111111111111;
			11'h4ef : dato = 32'b11111111111111111100010001100110;
			11'h4f0 : dato = 32'b01100110011001100110011001100110;
			11'h4f1 : dato = 32'b01100110011001100110011001100110;
			11'h4f2 : dato = 32'b01100110011001100110011001100110;
			11'h4f3 : dato = 32'b01100110011001100110011001100110;
			11'h4f4 : dato = 32'b01100110011001100110011001100110;
			11'h4f5 : dato = 32'b01100110011001100110011001100110;
			11'h4f6 : dato = 32'b01100110011001100110011001100110;
			11'h4f7 : dato = 32'b01100110011001100110011001100110;
			11'h4f8 : dato = 32'b01100110011001100110011001100110;
			11'h4f9 : dato = 32'b01100110011001100110011001100110;
			11'h4fa : dato = 32'b01100110011001100110011001100110;
			11'h4fb : dato = 32'b01100110011001100110011001100110;
			11'h4fc : dato = 32'b01100110011001100110110011110001;
			11'h4fd : dato = 32'b11111111111111111111111111111111;
			11'h4fe : dato = 32'b11111111111111111111111111111111;
			11'h4ff : dato = 32'b11111111111111111111111111111111;
			11'h500 : dato = 32'b11111111111111111111111111111111;
			11'h501 : dato = 32'b11111111111111111111111111111111;
			11'h502 : dato = 32'b11111111111111111111111111111111;
			11'h503 : dato = 32'b11111111111111111111110001111110;
			11'h504 : dato = 32'b01100110011001100110011001100110;
			11'h505 : dato = 32'b01100110011001100110011001100110;
			11'h506 : dato = 32'b01100110011001100110011001100110;
			11'h507 : dato = 32'b01100110011001100110011001100110;
			11'h508 : dato = 32'b01100110011001100110011001100110;
			11'h509 : dato = 32'b01100110011001100110011001100110;
			11'h50a : dato = 32'b01100110011001100110011001100110;
			11'h50b : dato = 32'b01100110011001100110011001100110;
			11'h50c : dato = 32'b01100110011001100110011001100110;
			11'h50d : dato = 32'b01100110011001100110011001100110;
			11'h50e : dato = 32'b01100110011001100110011001100110;
			11'h50f : dato = 32'b01100110011001100110011001100110;
			11'h510 : dato = 32'b01100110011001101010011111111111;
			11'h511 : dato = 32'b11111111111111111111111111111111;
			11'h512 : dato = 32'b11111111111111111111111111111111;
			11'h513 : dato = 32'b11111111111111111111111111111111;
			11'h514 : dato = 32'b11111111111111111111111111111111;
			11'h515 : dato = 32'b11111111111111111111111111111111;
			11'h516 : dato = 32'b11111111111111111111111111111111;
			11'h517 : dato = 32'b11111111111111111111111111011111;
			11'h518 : dato = 32'b01101010011001100110011001100110;
			11'h519 : dato = 32'b01100110011001100110011001100110;
			11'h51a : dato = 32'b01100110011001100110011001100110;
			11'h51b : dato = 32'b01100110011001100110011001100110;
			11'h51c : dato = 32'b01100110011001100110011001100110;
			11'h51d : dato = 32'b01100110011001100110011001100110;
			11'h51e : dato = 32'b01100110011001100110011001100110;
			11'h51f : dato = 32'b01100110011001100110011001100110;
			11'h520 : dato = 32'b01100110011001100110011001100110;
			11'h521 : dato = 32'b01100110011001100110011001100110;
			11'h522 : dato = 32'b01100110011001100110011001100110;
			11'h523 : dato = 32'b01100110011001100110011001100110;
			11'h524 : dato = 32'b01100110011011001110110111111111;
			11'h525 : dato = 32'b11111111111111111111111111111111;
			11'h526 : dato = 32'b11111111111111111111111111111111;
			11'h527 : dato = 32'b11111111111111111111111111111111;
			11'h528 : dato = 32'b11111111111111111111111111111111;
			11'h529 : dato = 32'b11111111111111111111111111111111;
			11'h52a : dato = 32'b11111111111111111111111111111111;
			11'h52b : dato = 32'b11111111111111111111111111111111;
			11'h52c : dato = 32'b10110010011001100110011001100110;
			11'h52d : dato = 32'b01100110011001100110011001100110;
			11'h52e : dato = 32'b01100110011001100110011001100110;
			11'h52f : dato = 32'b01100110011001100110011001100110;
			11'h530 : dato = 32'b01100110011001100110011001100110;
			11'h531 : dato = 32'b01100110011001100110011001100110;
			11'h532 : dato = 32'b01100110011001100110011001100110;
			11'h533 : dato = 32'b01100110011001100110011001100110;
			11'h534 : dato = 32'b01100110011001100110011001100110;
			11'h535 : dato = 32'b01100110011001100110011001100110;
			11'h536 : dato = 32'b01100110011001100110011001100110;
			11'h537 : dato = 32'b01100110011001100110011001100110;
			11'h538 : dato = 32'b01100110101110001111111111111111;
			11'h539 : dato = 32'b11111111111111111111111111111111;
			11'h53a : dato = 32'b11111111111111111111111111111111;
			11'h53b : dato = 32'b11111111111111111111111111111111;
			11'h53c : dato = 32'b11111111111111111111111111111111;
			11'h53d : dato = 32'b11111111111111111111111111111111;
			11'h53e : dato = 32'b11111111111111111111111111111111;
			11'h53f : dato = 32'b11111111111111111111111111111111;
			11'h540 : dato = 32'b11111100100000110110011001100110;
			11'h541 : dato = 32'b01100110011001100110011001100110;
			11'h542 : dato = 32'b01100110011001100110011001100110;
			11'h543 : dato = 32'b01100110011001100110011001100110;
			11'h544 : dato = 32'b01100110011001100110011001100110;
			11'h545 : dato = 32'b01100110011001100110011001100110;
			11'h546 : dato = 32'b01100110011001100110011001100110;
			11'h547 : dato = 32'b01100110011001100110011001100110;
			11'h548 : dato = 32'b01100110011001100110011001100110;
			11'h549 : dato = 32'b01100110011001100110011001100110;
			11'h54a : dato = 32'b01100110011001100110011001100110;
			11'h54b : dato = 32'b01100110011001100110011001100110;
			11'h54c : dato = 32'b10001110111111011111111111111111;
			11'h54d : dato = 32'b11111111111111111111111111111111;
			11'h54e : dato = 32'b11111111111111111111111111111111;
			11'h54f : dato = 32'b11111111111111111111111111111111;
			11'h550 : dato = 32'b11111111111111111111111111111111;
			11'h551 : dato = 32'b11111111111111111111111111111111;
			11'h552 : dato = 32'b11111111111111111111111111111111;
			11'h553 : dato = 32'b11111111111111111111111111111111;
			11'h554 : dato = 32'b11111111110111010110011001100110;
			11'h555 : dato = 32'b01100110011001100110011001100110;
			11'h556 : dato = 32'b01100110011001100110011001100110;
			11'h557 : dato = 32'b01100110011001100110011001100110;
			11'h558 : dato = 32'b01100110011001100110011001100110;
			11'h559 : dato = 32'b01100110011001100110011001100110;
			11'h55a : dato = 32'b01100110011001100110011001100110;
			11'h55b : dato = 32'b01100110011001100110011001100110;
			11'h55c : dato = 32'b01100110011001100110011001100110;
			11'h55d : dato = 32'b01100110011001100110011001100110;
			11'h55e : dato = 32'b01100110011001100110011001100110;
			11'h55f : dato = 32'b01100110011001100110011001110010;
			11'h560 : dato = 32'b11110100111111111111111111111111;
			11'h561 : dato = 32'b11111111111111111111111111111111;
			11'h562 : dato = 32'b11111111111111111111111111111111;
			11'h563 : dato = 32'b11111111111111111111111111111111;
			11'h564 : dato = 32'b11111111111111111111111111111111;
			11'h565 : dato = 32'b11111111111111111111111111111111;
			11'h566 : dato = 32'b11111111111111111111111111111111;
			11'h567 : dato = 32'b11111111111111111111111111111111;
			11'h568 : dato = 32'b11111111111111111010011001100110;
			11'h569 : dato = 32'b01100110011001100110011001100110;
			11'h56a : dato = 32'b01100110011001100110011001100110;
			11'h56b : dato = 32'b01100110011001100110011001100110;
			11'h56c : dato = 32'b01100110011001100110011001100110;
			11'h56d : dato = 32'b01100110011001100110011001100110;
			11'h56e : dato = 32'b01100110011001100110011001100110;
			11'h56f : dato = 32'b01100110011001100110011001100110;
			11'h570 : dato = 32'b01100110011001100110011001100110;
			11'h571 : dato = 32'b01100110011001100110011001100110;
			11'h572 : dato = 32'b01100110011001100110011001100110;
			11'h573 : dato = 32'b01100110011001100110011011001011;
			11'h574 : dato = 32'b11111111111111111111111111111111;
			11'h575 : dato = 32'b11111111111111111111111111111111;
			11'h576 : dato = 32'b11111111111111111111111111111111;
			11'h577 : dato = 32'b11111111111111111111111111111111;
			11'h578 : dato = 32'b11111111111111111111111111111111;
			11'h579 : dato = 32'b11111111111111111111111111111111;
			11'h57a : dato = 32'b11111111111111111111111111111111;
			11'h57b : dato = 32'b11111111111111111111111111111111;
			11'h57c : dato = 32'b11111111111111111111101110010000;
			11'h57d : dato = 32'b01100110011001100110011001100110;
			11'h57e : dato = 32'b01100110011001100110011001100110;
			11'h57f : dato = 32'b01100110011001100110011001100110;
			11'h580 : dato = 32'b01100110011001100110011001100110;
			11'h581 : dato = 32'b01100110011001100110011001100110;
			11'h582 : dato = 32'b01100110011001100110011001100110;
			11'h583 : dato = 32'b01100110011001100110011001100110;
			11'h584 : dato = 32'b01100110011001100110011001100110;
			11'h585 : dato = 32'b01100110011001100110011001100110;
			11'h586 : dato = 32'b01100110011001100110011001100110;
			11'h587 : dato = 32'b01100110011001101010100011111111;
			11'h588 : dato = 32'b11111111111111111111111111111111;
			11'h589 : dato = 32'b11111111111111111111111111111111;
			11'h58a : dato = 32'b11111111111111111111111111111111;
			11'h58b : dato = 32'b11111111111111111111111111111111;
			11'h58c : dato = 32'b11111111111111111111111111111111;
			11'h58d : dato = 32'b11111111111111111111111111111111;
			11'h58e : dato = 32'b11111111111111111111111111111111;
			11'h58f : dato = 32'b11111111111111111111111111111111;
			11'h590 : dato = 32'b11111111111111111111111111111011;
			11'h591 : dato = 32'b01111011011001100110011001100110;
			11'h592 : dato = 32'b01100110011001100110011001100110;
			11'h593 : dato = 32'b01100110011001100110011001100110;
			11'h594 : dato = 32'b01100110011001100110011001100110;
			11'h595 : dato = 32'b01100110011001100110011001100110;
			11'h596 : dato = 32'b01100110011001100110011001100110;
			11'h597 : dato = 32'b01100110011001100110011001100110;
			11'h598 : dato = 32'b01100110011001100110011001100110;
			11'h599 : dato = 32'b01100110011001100110011001100110;
			11'h59a : dato = 32'b01100110011001100110011001100110;
			11'h59b : dato = 32'b01100110100011111111110011111111;
			11'h59c : dato = 32'b11111111111111111111111111111111;
			11'h59d : dato = 32'b11111111111111111111111111111111;
			11'h59e : dato = 32'b11111111111111111111111111111111;
			11'h59f : dato = 32'b11111111111111111111111111111111;
			11'h5a0 : dato = 32'b11111111111111111111111111111111;
			11'h5a1 : dato = 32'b11111111111111111111111111111111;
			11'h5a2 : dato = 32'b11111111111111111111111111111111;
			11'h5a3 : dato = 32'b11111111111111111111111111111111;
			11'h5a4 : dato = 32'b11111111111111111111111111111111;
			11'h5a5 : dato = 32'b11110011100000100110011001100110;
			11'h5a6 : dato = 32'b01100110011001100110011001100110;
			11'h5a7 : dato = 32'b01100110011001100110011001100110;
			11'h5a8 : dato = 32'b01100110011001100110011001100110;
			11'h5a9 : dato = 32'b01100110011001100110011001100110;
			11'h5aa : dato = 32'b01100110011001100110011001100110;
			11'h5ab : dato = 32'b01100110011001100110011001100110;
			11'h5ac : dato = 32'b01100110011001100110011001100110;
			11'h5ad : dato = 32'b01100110011001100110011001100110;
			11'h5ae : dato = 32'b01100110011001100110011001100110;
			11'h5af : dato = 32'b10000100111101111111111111111111;
			11'h5b0 : dato = 32'b11111111111111111111111111111111;
			11'h5b1 : dato = 32'b11111111111111111111111111111111;
			11'h5b2 : dato = 32'b11111111111111111111111111111111;
			11'h5b3 : dato = 32'b11111111111111111111111111111111;
			11'h5b4 : dato = 32'b11111111111111111111111111111111;
			11'h5b5 : dato = 32'b11111111111111111111111111111111;
			11'h5b6 : dato = 32'b11111111111111111111111111111111;
			11'h5b7 : dato = 32'b11111111111111111111111111111111;
			11'h5b8 : dato = 32'b11111111111111111111111111111111;
			11'h5b9 : dato = 32'b11111111111011110111001101100110;
			11'h5ba : dato = 32'b01100110011001100110011001100110;
			11'h5bb : dato = 32'b01100110011001100110011001100110;
			11'h5bc : dato = 32'b01100110011001100110011001100110;
			11'h5bd : dato = 32'b01100110011001100110011010000000;
			11'h5be : dato = 32'b10001110100010110111001101100110;
			11'h5bf : dato = 32'b01100110011001100110011001100110;
			11'h5c0 : dato = 32'b01100110011001100110011001100110;
			11'h5c1 : dato = 32'b01100110011001100110011001100110;
			11'h5c2 : dato = 32'b01100110011001100110011001111011;
			11'h5c3 : dato = 32'b11101111111111111111111111111111;
			11'h5c4 : dato = 32'b11111111111111111111111111111111;
			11'h5c5 : dato = 32'b11111111111111111111111111111111;
			11'h5c6 : dato = 32'b11111111111111111111111111111111;
			11'h5c7 : dato = 32'b11111111111111111111111111111111;
			11'h5c8 : dato = 32'b11111111111111111111111111111111;
			11'h5c9 : dato = 32'b11111111111111111111111111111111;
			11'h5ca : dato = 32'b11111111111111111111111111111111;
			11'h5cb : dato = 32'b11111111111111111111111111111111;
			11'h5cc : dato = 32'b11111111111111111111111111111111;
			11'h5cd : dato = 32'b11111111111111111110010001111011;
			11'h5ce : dato = 32'b01100110011001100110011001100110;
			11'h5cf : dato = 32'b01100110011001100110011001100110;
			11'h5d0 : dato = 32'b01100110011001100110011010000000;
			11'h5d1 : dato = 32'b10101110110101011111010111111111;
			11'h5d2 : dato = 32'b11111111111111111111111111110000;
			11'h5d3 : dato = 32'b11001100101000110111111001100110;
			11'h5d4 : dato = 32'b01100110011001100110011001100110;
			11'h5d5 : dato = 32'b01100110011001100110011001100110;
			11'h5d6 : dato = 32'b01100110011001101001010011110100;
			11'h5d7 : dato = 32'b11111111111111111111111111111111;
			11'h5d8 : dato = 32'b11111111111111111111111111111111;
			11'h5d9 : dato = 32'b11111111111111111111111111111111;
			11'h5da : dato = 32'b11111111111111111111111111111111;
			11'h5db : dato = 32'b11111111111111111111111111111111;
			11'h5dc : dato = 32'b11111111111111111111111111111111;
			11'h5dd : dato = 32'b11111111111111111111111111111111;
			11'h5de : dato = 32'b11111111111111111111111111111111;
			11'h5df : dato = 32'b11111111111111111111111111111111;
			11'h5e0 : dato = 32'b11111111111111111111111111111111;
			11'h5e1 : dato = 32'b11111111111111111111111111110111;
			11'h5e2 : dato = 32'b10110101011101000110011001100110;
			11'h5e3 : dato = 32'b01100110011001100110011001101100;
			11'h5e4 : dato = 32'b10010100101110111110010111111111;
			11'h5e5 : dato = 32'b11111111111111111111111111111111;
			11'h5e6 : dato = 32'b11111111111111111111111111111111;
			11'h5e7 : dato = 32'b11111111111111111111111111101100;
			11'h5e8 : dato = 32'b10111001100010000110100001100110;
			11'h5e9 : dato = 32'b01100110011001100110011001100110;
			11'h5ea : dato = 32'b01110001110000001111111011111111;
			11'h5eb : dato = 32'b11111111111111111111111111111111;
			11'h5ec : dato = 32'b11111111111111111111111111111111;
			11'h5ed : dato = 32'b11111111111111111111111111111111;
			11'h5ee : dato = 32'b11111111111111111111111111111111;
			11'h5ef : dato = 32'b11111111111111111111111111111111;
			11'h5f0 : dato = 32'b11111111111111111111111111111111;
			11'h5f1 : dato = 32'b11111111111111111111111111111111;
			11'h5f2 : dato = 32'b11111111111111111111111111111111;
			11'h5f3 : dato = 32'b11111111111111111111111111111111;
			11'h5f4 : dato = 32'b11111111111111111111111111111111;
			11'h5f5 : dato = 32'b11111111111111111111111111111111;
			11'h5f6 : dato = 32'b11111111111110111101000010101101;
			11'h5f7 : dato = 32'b10100010101100101101011111111011;
			11'h5f8 : dato = 32'b11111111111111111111111111111111;
			11'h5f9 : dato = 32'b11111111111111111111111111111111;
			11'h5fa : dato = 32'b11111111111111111111111111111111;
			11'h5fb : dato = 32'b11111111111111111111111111111111;
			11'h5fc : dato = 32'b11111111111111111111011011011000;
			11'h5fd : dato = 32'b11000001101100111011011011010000;
			11'h5fe : dato = 32'b11111001111111111111111111111111;
			11'h5ff : dato = 32'b11111111111111111111111111111111;
			11'h600 : dato = 32'b11111111111111111111111111111111;
			11'h601 : dato = 32'b11111111111111111111111111111111;
			11'h602 : dato = 32'b11111111111111111111111111111111;
			11'h603 : dato = 32'b11111111111111111111111111111111;
			11'h604 : dato = 32'b11111111111111111111111111111111;
			11'h605 : dato = 32'b11111111111111111111111111111111;
			11'h606 : dato = 32'b11111111111111111111111111111111;
			11'h607 : dato = 32'b11111111111111111111111111111111;
			11'h608 : dato = 32'b11111111111111111111111111111111;
			11'h609 : dato = 32'b11111111111111111111111111111111;
			11'h60a : dato = 32'b11111111111111111111111111111111;
			11'h60b : dato = 32'b11111111111111111111111111111111;
			11'h60c : dato = 32'b11111111111111111111111111111111;
			11'h60d : dato = 32'b11111111111111111111111111111111;
			11'h60e : dato = 32'b11111111111111111111111111111111;
			11'h60f : dato = 32'b11111111111111111111111111111111;
			11'h610 : dato = 32'b11111111111111111111111111111111;
			11'h611 : dato = 32'b11111111111111111111111111111111;
			11'h612 : dato = 32'b11111111111111111111111111111111;
			11'h613 : dato = 32'b11111111111111111111111111111111;
			11'h614 : dato = 32'b11111111111111111111111111111111;
			11'h615 : dato = 32'b11111111111111111111111111111111;
			11'h616 : dato = 32'b11111111111111111111111111111111;
			11'h617 : dato = 32'b11111111111111111111111111111111;
			11'h618 : dato = 32'b11111111111111111111111111111111;
			11'h619 : dato = 32'b11111111111111111111111111111111;
			11'h61a : dato = 32'b11111111111111111111111111111111;
			11'h61b : dato = 32'b11111111111111111111111111111111;
			11'h61c : dato = 32'b11111111111111111111111111111111;
			11'h61d : dato = 32'b11111111111111111111111111111111;
			11'h61e : dato = 32'b11111111111111111111111111111111;
			11'h61f : dato = 32'b11111111111111111111111111111111;
			11'h620 : dato = 32'b11111111111111111111111111111111;
			11'h621 : dato = 32'b11111111111111111111111111111111;
			11'h622 : dato = 32'b11111111111111111111111111111111;
			11'h623 : dato = 32'b11111111111111111111111111111111;
			11'h624 : dato = 32'b11111111111111111111111111111111;
			11'h625 : dato = 32'b11111111111111111111111111111111;
			11'h626 : dato = 32'b11111111111111111111111111111111;
			11'h627 : dato = 32'b11111111111111111111111111111111;
			11'h628 : dato = 32'b11111111111111111111111111111111;
			11'h629 : dato = 32'b11111111111111111111111111111111;
			11'h62a : dato = 32'b11111111111111111111111111111111;
			11'h62b : dato = 32'b11111111111111111111111111111111;
			11'h62c : dato = 32'b11111111111111111111111111111111;
			11'h62d : dato = 32'b11111111111111111111111111111111;
			11'h62e : dato = 32'b11111111111111111111111111111111;
			11'h62f : dato = 32'b11111111111111111111111111111111;
			11'h630 : dato = 32'b11111111111111111111111111111111;
			11'h631 : dato = 32'b11111111111111111111111111111111;
			11'h632 : dato = 32'b11111111111111111111111111111111;
			11'h633 : dato = 32'b11111111111111111111111111111111;
			11'h634 : dato = 32'b11111111111111111111111111111111;
			11'h635 : dato = 32'b11111111111111111111111111111111;
			11'h636 : dato = 32'b11111111111111111111111111111111;
			11'h637 : dato = 32'b11111111111111111111111111111111;
			11'h638 : dato = 32'b11111111111111111111111111111111;
			11'h639 : dato = 32'b11111111111111111111111111111111;
			11'h63a : dato = 32'b11111111111111111111111111111111;
			11'h63b : dato = 32'b11111111111111111111111111111111;
			11'h63c : dato = 32'b11111111111111111111111111111111;
			11'h63d : dato = 32'b11111111111111111111111111111111;
			11'h63e : dato = 32'b11111111111111111111111111111111;
			11'h63f : dato = 32'b11111111111111111111111111111111;
			default: dato = 32'b1;
		endcase

endmodule