logic [1:0] sprite [0:123][0:99] = 
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}}
'{'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}}
'{'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}}
'{'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b11}'{2'b11}'{2'b11}'{2'b11}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b10}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
'{'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b01}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}'{2'b00}}
;